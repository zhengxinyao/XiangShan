module PayloadArray(
  input         clock,
  input  [15:0] io_read_0_addr,
  output [9:0]  io_read_0_data_cf_foldpc,
  output        io_read_0_data_cf_trigger_backendEn_0,
  output        io_read_0_data_cf_trigger_backendEn_1,
  output        io_read_0_data_cf_pd_isRVC,
  output [1:0]  io_read_0_data_cf_pd_brType,
  output        io_read_0_data_cf_pd_isCall,
  output        io_read_0_data_cf_pd_isRet,
  output        io_read_0_data_cf_pred_taken,
  output        io_read_0_data_cf_storeSetHit,
  output        io_read_0_data_cf_waitForRobIdx_flag,
  output [4:0]  io_read_0_data_cf_waitForRobIdx_value,
  output        io_read_0_data_cf_loadWaitBit,
  output        io_read_0_data_cf_loadWaitStrict,
  output [4:0]  io_read_0_data_cf_ssid,
  output        io_read_0_data_cf_ftqPtr_flag,
  output [2:0]  io_read_0_data_cf_ftqPtr_value,
  output [2:0]  io_read_0_data_cf_ftqOffset,
  output [3:0]  io_read_0_data_ctrl_fuType,
  output [6:0]  io_read_0_data_ctrl_fuOpType,
  output        io_read_0_data_ctrl_rfWen,
  output        io_read_0_data_ctrl_fpWen,
  output [19:0] io_read_0_data_ctrl_imm,
  output [5:0]  io_read_0_data_pdest,
  output        io_read_0_data_robIdx_flag,
  output [4:0]  io_read_0_data_robIdx_value,
  output        io_read_0_data_lqIdx_flag,
  output [3:0]  io_read_0_data_lqIdx_value,
  output        io_read_0_data_sqIdx_flag,
  output [3:0]  io_read_0_data_sqIdx_value,
  input  [15:0] io_read_1_addr,
  output [9:0]  io_read_1_data_cf_foldpc,
  output        io_read_1_data_cf_trigger_backendEn_0,
  output        io_read_1_data_cf_trigger_backendEn_1,
  output        io_read_1_data_cf_pd_isRVC,
  output [1:0]  io_read_1_data_cf_pd_brType,
  output        io_read_1_data_cf_pd_isCall,
  output        io_read_1_data_cf_pd_isRet,
  output        io_read_1_data_cf_pred_taken,
  output        io_read_1_data_cf_storeSetHit,
  output        io_read_1_data_cf_waitForRobIdx_flag,
  output [4:0]  io_read_1_data_cf_waitForRobIdx_value,
  output        io_read_1_data_cf_loadWaitBit,
  output        io_read_1_data_cf_loadWaitStrict,
  output [4:0]  io_read_1_data_cf_ssid,
  output        io_read_1_data_cf_ftqPtr_flag,
  output [2:0]  io_read_1_data_cf_ftqPtr_value,
  output [2:0]  io_read_1_data_cf_ftqOffset,
  output [3:0]  io_read_1_data_ctrl_fuType,
  output [6:0]  io_read_1_data_ctrl_fuOpType,
  output        io_read_1_data_ctrl_rfWen,
  output        io_read_1_data_ctrl_fpWen,
  output [19:0] io_read_1_data_ctrl_imm,
  output [5:0]  io_read_1_data_pdest,
  output        io_read_1_data_robIdx_flag,
  output [4:0]  io_read_1_data_robIdx_value,
  output        io_read_1_data_lqIdx_flag,
  output [3:0]  io_read_1_data_lqIdx_value,
  output        io_read_1_data_sqIdx_flag,
  output [3:0]  io_read_1_data_sqIdx_value,
  input  [15:0] io_read_2_addr,
  output [9:0]  io_read_2_data_cf_foldpc,
  output        io_read_2_data_cf_trigger_backendEn_0,
  output        io_read_2_data_cf_trigger_backendEn_1,
  output        io_read_2_data_cf_pd_isRVC,
  output [1:0]  io_read_2_data_cf_pd_brType,
  output        io_read_2_data_cf_pd_isCall,
  output        io_read_2_data_cf_pd_isRet,
  output        io_read_2_data_cf_pred_taken,
  output        io_read_2_data_cf_storeSetHit,
  output        io_read_2_data_cf_waitForRobIdx_flag,
  output [4:0]  io_read_2_data_cf_waitForRobIdx_value,
  output        io_read_2_data_cf_loadWaitBit,
  output        io_read_2_data_cf_loadWaitStrict,
  output [4:0]  io_read_2_data_cf_ssid,
  output        io_read_2_data_cf_ftqPtr_flag,
  output [2:0]  io_read_2_data_cf_ftqPtr_value,
  output [2:0]  io_read_2_data_cf_ftqOffset,
  output [3:0]  io_read_2_data_ctrl_fuType,
  output [6:0]  io_read_2_data_ctrl_fuOpType,
  output        io_read_2_data_ctrl_rfWen,
  output        io_read_2_data_ctrl_fpWen,
  output [19:0] io_read_2_data_ctrl_imm,
  output [5:0]  io_read_2_data_pdest,
  output        io_read_2_data_robIdx_flag,
  output [4:0]  io_read_2_data_robIdx_value,
  output        io_read_2_data_lqIdx_flag,
  output [3:0]  io_read_2_data_lqIdx_value,
  output        io_read_2_data_sqIdx_flag,
  output [3:0]  io_read_2_data_sqIdx_value,
  input         io_write_0_enable,
  input  [15:0] io_write_0_addr,
  input  [9:0]  io_write_0_data_cf_foldpc,
  input         io_write_0_data_cf_trigger_backendEn_0,
  input         io_write_0_data_cf_trigger_backendEn_1,
  input         io_write_0_data_cf_pd_isRVC,
  input  [1:0]  io_write_0_data_cf_pd_brType,
  input         io_write_0_data_cf_pd_isCall,
  input         io_write_0_data_cf_pd_isRet,
  input         io_write_0_data_cf_pred_taken,
  input         io_write_0_data_cf_storeSetHit,
  input         io_write_0_data_cf_waitForRobIdx_flag,
  input  [4:0]  io_write_0_data_cf_waitForRobIdx_value,
  input         io_write_0_data_cf_loadWaitBit,
  input         io_write_0_data_cf_loadWaitStrict,
  input  [4:0]  io_write_0_data_cf_ssid,
  input         io_write_0_data_cf_ftqPtr_flag,
  input  [2:0]  io_write_0_data_cf_ftqPtr_value,
  input  [2:0]  io_write_0_data_cf_ftqOffset,
  input  [3:0]  io_write_0_data_ctrl_fuType,
  input  [6:0]  io_write_0_data_ctrl_fuOpType,
  input         io_write_0_data_ctrl_rfWen,
  input         io_write_0_data_ctrl_fpWen,
  input  [19:0] io_write_0_data_ctrl_imm,
  input  [5:0]  io_write_0_data_pdest,
  input         io_write_0_data_robIdx_flag,
  input  [4:0]  io_write_0_data_robIdx_value,
  input         io_write_0_data_lqIdx_flag,
  input  [3:0]  io_write_0_data_lqIdx_value,
  input         io_write_0_data_sqIdx_flag,
  input  [3:0]  io_write_0_data_sqIdx_value,
  input         io_write_1_enable,
  input  [15:0] io_write_1_addr,
  input  [9:0]  io_write_1_data_cf_foldpc,
  input         io_write_1_data_cf_trigger_backendEn_0,
  input         io_write_1_data_cf_trigger_backendEn_1,
  input         io_write_1_data_cf_pd_isRVC,
  input  [1:0]  io_write_1_data_cf_pd_brType,
  input         io_write_1_data_cf_pd_isCall,
  input         io_write_1_data_cf_pd_isRet,
  input         io_write_1_data_cf_pred_taken,
  input         io_write_1_data_cf_storeSetHit,
  input         io_write_1_data_cf_waitForRobIdx_flag,
  input  [4:0]  io_write_1_data_cf_waitForRobIdx_value,
  input         io_write_1_data_cf_loadWaitBit,
  input         io_write_1_data_cf_loadWaitStrict,
  input  [4:0]  io_write_1_data_cf_ssid,
  input         io_write_1_data_cf_ftqPtr_flag,
  input  [2:0]  io_write_1_data_cf_ftqPtr_value,
  input  [2:0]  io_write_1_data_cf_ftqOffset,
  input  [3:0]  io_write_1_data_ctrl_fuType,
  input  [6:0]  io_write_1_data_ctrl_fuOpType,
  input         io_write_1_data_ctrl_rfWen,
  input         io_write_1_data_ctrl_fpWen,
  input  [19:0] io_write_1_data_ctrl_imm,
  input  [5:0]  io_write_1_data_pdest,
  input         io_write_1_data_robIdx_flag,
  input  [4:0]  io_write_1_data_robIdx_value,
  input         io_write_1_data_lqIdx_flag,
  input  [3:0]  io_write_1_data_lqIdx_value,
  input         io_write_1_data_sqIdx_flag,
  input  [3:0]  io_write_1_data_sqIdx_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] payload_0_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_0_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_0_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_0_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_0_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_0_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_0_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_0_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_0_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_0_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_0_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_0_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_0_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_0_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_0_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_0_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_1_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_1_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_1_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_1_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_1_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_1_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_1_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_1_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_1_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_1_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_1_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_1_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_1_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_1_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_1_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_1_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_2_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_2_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_2_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_2_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_2_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_2_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_2_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_2_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_2_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_2_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_2_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_2_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_2_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_2_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_2_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_2_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_3_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_3_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_3_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_3_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_3_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_3_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_3_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_3_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_3_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_3_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_3_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_3_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_3_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_3_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_3_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_3_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_4_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_4_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_4_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_4_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_4_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_4_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_4_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_4_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_4_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_4_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_4_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_4_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_4_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_4_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_4_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_4_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_5_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_5_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_5_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_5_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_5_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_5_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_5_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_5_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_5_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_5_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_5_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_5_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_5_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_5_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_5_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_5_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_6_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_6_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_6_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_6_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_6_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_6_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_6_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_6_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_6_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_6_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_6_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_6_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_6_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_6_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_6_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_6_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_7_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_7_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_7_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_7_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_7_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_7_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_7_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_7_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_7_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_7_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_7_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_7_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_7_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_7_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_7_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_7_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_8_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_8_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_8_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_8_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_8_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_8_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_8_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_8_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_8_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_8_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_8_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_8_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_8_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_8_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_8_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_8_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_8_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_8_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_8_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_9_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_9_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_9_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_9_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_9_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_9_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_9_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_9_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_9_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_9_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_9_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_9_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_9_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_9_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_9_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_9_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_9_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_9_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_9_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_10_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_10_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_10_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_10_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_10_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_10_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_10_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_10_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_10_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_10_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_10_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_10_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_10_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_10_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_10_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_10_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_10_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_10_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_10_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_11_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_11_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_11_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_11_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_11_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_11_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_11_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_11_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_11_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_11_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_11_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_11_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_11_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_11_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_11_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_11_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_11_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_11_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_11_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_12_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_12_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_12_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_12_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_12_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_12_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_12_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_12_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_12_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_12_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_12_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_12_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_12_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_12_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_12_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_12_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_12_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_12_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_12_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_13_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_13_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_13_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_13_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_13_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_13_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_13_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_13_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_13_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_13_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_13_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_13_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_13_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_13_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_13_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_13_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_13_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_13_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_13_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_14_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_14_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_14_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_14_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_14_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_14_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_14_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_14_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_14_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_14_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_14_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_14_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_14_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_14_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_14_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_14_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_14_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_14_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_14_sqIdx_value; // @[PayloadArray.scala 45:20]
  reg [9:0] payload_15_cf_foldpc; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_trigger_backendEn_0; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_trigger_backendEn_1; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_15_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_storeSetHit; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_waitForRobIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_15_cf_waitForRobIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_loadWaitBit; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_loadWaitStrict; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_15_cf_ssid; // @[PayloadArray.scala 45:20]
  reg  payload_15_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_15_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_15_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_15_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_15_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_15_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_15_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_15_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_15_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_15_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_15_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_15_lqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_15_lqIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_15_sqIdx_flag; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_15_sqIdx_value; // @[PayloadArray.scala 45:20]
  wire [3:0] _io_read_0_data_T_357 = io_read_0_addr[0] ? payload_0_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_358 = io_read_0_addr[1] ? payload_1_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_359 = io_read_0_addr[2] ? payload_2_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_360 = io_read_0_addr[3] ? payload_3_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_361 = io_read_0_addr[4] ? payload_4_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_362 = io_read_0_addr[5] ? payload_5_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_363 = io_read_0_addr[6] ? payload_6_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_364 = io_read_0_addr[7] ? payload_7_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_365 = io_read_0_addr[8] ? payload_8_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_366 = io_read_0_addr[9] ? payload_9_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_367 = io_read_0_addr[10] ? payload_10_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_368 = io_read_0_addr[11] ? payload_11_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_369 = io_read_0_addr[12] ? payload_12_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_370 = io_read_0_addr[13] ? payload_13_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_371 = io_read_0_addr[14] ? payload_14_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_372 = io_read_0_addr[15] ? payload_15_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_373 = _io_read_0_data_T_357 | _io_read_0_data_T_358; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_374 = _io_read_0_data_T_373 | _io_read_0_data_T_359; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_375 = _io_read_0_data_T_374 | _io_read_0_data_T_360; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_376 = _io_read_0_data_T_375 | _io_read_0_data_T_361; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_377 = _io_read_0_data_T_376 | _io_read_0_data_T_362; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_378 = _io_read_0_data_T_377 | _io_read_0_data_T_363; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_379 = _io_read_0_data_T_378 | _io_read_0_data_T_364; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_380 = _io_read_0_data_T_379 | _io_read_0_data_T_365; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_381 = _io_read_0_data_T_380 | _io_read_0_data_T_366; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_382 = _io_read_0_data_T_381 | _io_read_0_data_T_367; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_383 = _io_read_0_data_T_382 | _io_read_0_data_T_368; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_384 = _io_read_0_data_T_383 | _io_read_0_data_T_369; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_385 = _io_read_0_data_T_384 | _io_read_0_data_T_370; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_386 = _io_read_0_data_T_385 | _io_read_0_data_T_371; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_403 = io_read_0_addr[15] & payload_15_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_419 = io_read_0_addr[0] ? payload_0_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_420 = io_read_0_addr[1] ? payload_1_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_421 = io_read_0_addr[2] ? payload_2_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_422 = io_read_0_addr[3] ? payload_3_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_423 = io_read_0_addr[4] ? payload_4_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_424 = io_read_0_addr[5] ? payload_5_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_425 = io_read_0_addr[6] ? payload_6_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_426 = io_read_0_addr[7] ? payload_7_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_427 = io_read_0_addr[8] ? payload_8_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_428 = io_read_0_addr[9] ? payload_9_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_429 = io_read_0_addr[10] ? payload_10_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_430 = io_read_0_addr[11] ? payload_11_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_431 = io_read_0_addr[12] ? payload_12_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_432 = io_read_0_addr[13] ? payload_13_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_433 = io_read_0_addr[14] ? payload_14_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_434 = io_read_0_addr[15] ? payload_15_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_435 = _io_read_0_data_T_419 | _io_read_0_data_T_420; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_436 = _io_read_0_data_T_435 | _io_read_0_data_T_421; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_437 = _io_read_0_data_T_436 | _io_read_0_data_T_422; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_438 = _io_read_0_data_T_437 | _io_read_0_data_T_423; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_439 = _io_read_0_data_T_438 | _io_read_0_data_T_424; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_440 = _io_read_0_data_T_439 | _io_read_0_data_T_425; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_441 = _io_read_0_data_T_440 | _io_read_0_data_T_426; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_442 = _io_read_0_data_T_441 | _io_read_0_data_T_427; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_443 = _io_read_0_data_T_442 | _io_read_0_data_T_428; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_444 = _io_read_0_data_T_443 | _io_read_0_data_T_429; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_445 = _io_read_0_data_T_444 | _io_read_0_data_T_430; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_446 = _io_read_0_data_T_445 | _io_read_0_data_T_431; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_447 = _io_read_0_data_T_446 | _io_read_0_data_T_432; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_448 = _io_read_0_data_T_447 | _io_read_0_data_T_433; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_465 = io_read_0_addr[15] & payload_15_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_481 = io_read_0_addr[0] ? payload_0_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_482 = io_read_0_addr[1] ? payload_1_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_483 = io_read_0_addr[2] ? payload_2_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_484 = io_read_0_addr[3] ? payload_3_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_485 = io_read_0_addr[4] ? payload_4_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_486 = io_read_0_addr[5] ? payload_5_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_487 = io_read_0_addr[6] ? payload_6_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_488 = io_read_0_addr[7] ? payload_7_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_489 = io_read_0_addr[8] ? payload_8_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_490 = io_read_0_addr[9] ? payload_9_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_491 = io_read_0_addr[10] ? payload_10_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_492 = io_read_0_addr[11] ? payload_11_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_493 = io_read_0_addr[12] ? payload_12_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_494 = io_read_0_addr[13] ? payload_13_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_495 = io_read_0_addr[14] ? payload_14_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_496 = io_read_0_addr[15] ? payload_15_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_497 = _io_read_0_data_T_481 | _io_read_0_data_T_482; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_498 = _io_read_0_data_T_497 | _io_read_0_data_T_483; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_499 = _io_read_0_data_T_498 | _io_read_0_data_T_484; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_500 = _io_read_0_data_T_499 | _io_read_0_data_T_485; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_501 = _io_read_0_data_T_500 | _io_read_0_data_T_486; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_502 = _io_read_0_data_T_501 | _io_read_0_data_T_487; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_503 = _io_read_0_data_T_502 | _io_read_0_data_T_488; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_504 = _io_read_0_data_T_503 | _io_read_0_data_T_489; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_505 = _io_read_0_data_T_504 | _io_read_0_data_T_490; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_506 = _io_read_0_data_T_505 | _io_read_0_data_T_491; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_507 = _io_read_0_data_T_506 | _io_read_0_data_T_492; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_508 = _io_read_0_data_T_507 | _io_read_0_data_T_493; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_509 = _io_read_0_data_T_508 | _io_read_0_data_T_494; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_510 = _io_read_0_data_T_509 | _io_read_0_data_T_495; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_527 = io_read_0_addr[15] & payload_15_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_574 = io_read_0_addr[0] ? payload_0_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_575 = io_read_0_addr[1] ? payload_1_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_576 = io_read_0_addr[2] ? payload_2_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_577 = io_read_0_addr[3] ? payload_3_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_578 = io_read_0_addr[4] ? payload_4_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_579 = io_read_0_addr[5] ? payload_5_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_580 = io_read_0_addr[6] ? payload_6_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_581 = io_read_0_addr[7] ? payload_7_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_582 = io_read_0_addr[8] ? payload_8_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_583 = io_read_0_addr[9] ? payload_9_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_584 = io_read_0_addr[10] ? payload_10_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_585 = io_read_0_addr[11] ? payload_11_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_586 = io_read_0_addr[12] ? payload_12_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_587 = io_read_0_addr[13] ? payload_13_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_588 = io_read_0_addr[14] ? payload_14_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_589 = io_read_0_addr[15] ? payload_15_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_590 = _io_read_0_data_T_574 | _io_read_0_data_T_575; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_591 = _io_read_0_data_T_590 | _io_read_0_data_T_576; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_592 = _io_read_0_data_T_591 | _io_read_0_data_T_577; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_593 = _io_read_0_data_T_592 | _io_read_0_data_T_578; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_594 = _io_read_0_data_T_593 | _io_read_0_data_T_579; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_595 = _io_read_0_data_T_594 | _io_read_0_data_T_580; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_596 = _io_read_0_data_T_595 | _io_read_0_data_T_581; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_597 = _io_read_0_data_T_596 | _io_read_0_data_T_582; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_598 = _io_read_0_data_T_597 | _io_read_0_data_T_583; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_599 = _io_read_0_data_T_598 | _io_read_0_data_T_584; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_600 = _io_read_0_data_T_599 | _io_read_0_data_T_585; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_601 = _io_read_0_data_T_600 | _io_read_0_data_T_586; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_602 = _io_read_0_data_T_601 | _io_read_0_data_T_587; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_603 = _io_read_0_data_T_602 | _io_read_0_data_T_588; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1349 = io_read_0_addr[0] ? payload_0_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1350 = io_read_0_addr[1] ? payload_1_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1351 = io_read_0_addr[2] ? payload_2_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1352 = io_read_0_addr[3] ? payload_3_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1353 = io_read_0_addr[4] ? payload_4_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1354 = io_read_0_addr[5] ? payload_5_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1355 = io_read_0_addr[6] ? payload_6_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1356 = io_read_0_addr[7] ? payload_7_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1357 = io_read_0_addr[8] ? payload_8_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1358 = io_read_0_addr[9] ? payload_9_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1359 = io_read_0_addr[10] ? payload_10_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1360 = io_read_0_addr[11] ? payload_11_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1361 = io_read_0_addr[12] ? payload_12_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1362 = io_read_0_addr[13] ? payload_13_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1363 = io_read_0_addr[14] ? payload_14_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1364 = io_read_0_addr[15] ? payload_15_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1365 = _io_read_0_data_T_1349 | _io_read_0_data_T_1350; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1366 = _io_read_0_data_T_1365 | _io_read_0_data_T_1351; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1367 = _io_read_0_data_T_1366 | _io_read_0_data_T_1352; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1368 = _io_read_0_data_T_1367 | _io_read_0_data_T_1353; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1369 = _io_read_0_data_T_1368 | _io_read_0_data_T_1354; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1370 = _io_read_0_data_T_1369 | _io_read_0_data_T_1355; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1371 = _io_read_0_data_T_1370 | _io_read_0_data_T_1356; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1372 = _io_read_0_data_T_1371 | _io_read_0_data_T_1357; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1373 = _io_read_0_data_T_1372 | _io_read_0_data_T_1358; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1374 = _io_read_0_data_T_1373 | _io_read_0_data_T_1359; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1375 = _io_read_0_data_T_1374 | _io_read_0_data_T_1360; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1376 = _io_read_0_data_T_1375 | _io_read_0_data_T_1361; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1377 = _io_read_0_data_T_1376 | _io_read_0_data_T_1362; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_1378 = _io_read_0_data_T_1377 | _io_read_0_data_T_1363; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_1550 = io_read_0_addr[15] & payload_15_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_1581 = io_read_0_addr[15] & payload_15_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1597 = io_read_0_addr[0] ? payload_0_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1598 = io_read_0_addr[1] ? payload_1_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1599 = io_read_0_addr[2] ? payload_2_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1600 = io_read_0_addr[3] ? payload_3_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1601 = io_read_0_addr[4] ? payload_4_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1602 = io_read_0_addr[5] ? payload_5_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1603 = io_read_0_addr[6] ? payload_6_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1604 = io_read_0_addr[7] ? payload_7_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1605 = io_read_0_addr[8] ? payload_8_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1606 = io_read_0_addr[9] ? payload_9_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1607 = io_read_0_addr[10] ? payload_10_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1608 = io_read_0_addr[11] ? payload_11_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1609 = io_read_0_addr[12] ? payload_12_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1610 = io_read_0_addr[13] ? payload_13_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1611 = io_read_0_addr[14] ? payload_14_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1612 = io_read_0_addr[15] ? payload_15_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1613 = _io_read_0_data_T_1597 | _io_read_0_data_T_1598; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1614 = _io_read_0_data_T_1613 | _io_read_0_data_T_1599; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1615 = _io_read_0_data_T_1614 | _io_read_0_data_T_1600; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1616 = _io_read_0_data_T_1615 | _io_read_0_data_T_1601; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1617 = _io_read_0_data_T_1616 | _io_read_0_data_T_1602; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1618 = _io_read_0_data_T_1617 | _io_read_0_data_T_1603; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1619 = _io_read_0_data_T_1618 | _io_read_0_data_T_1604; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1620 = _io_read_0_data_T_1619 | _io_read_0_data_T_1605; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1621 = _io_read_0_data_T_1620 | _io_read_0_data_T_1606; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1622 = _io_read_0_data_T_1621 | _io_read_0_data_T_1607; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1623 = _io_read_0_data_T_1622 | _io_read_0_data_T_1608; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1624 = _io_read_0_data_T_1623 | _io_read_0_data_T_1609; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1625 = _io_read_0_data_T_1624 | _io_read_0_data_T_1610; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_1626 = _io_read_0_data_T_1625 | _io_read_0_data_T_1611; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1628 = io_read_0_addr[0] ? payload_0_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1629 = io_read_0_addr[1] ? payload_1_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1630 = io_read_0_addr[2] ? payload_2_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1631 = io_read_0_addr[3] ? payload_3_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1632 = io_read_0_addr[4] ? payload_4_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1633 = io_read_0_addr[5] ? payload_5_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1634 = io_read_0_addr[6] ? payload_6_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1635 = io_read_0_addr[7] ? payload_7_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1636 = io_read_0_addr[8] ? payload_8_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1637 = io_read_0_addr[9] ? payload_9_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1638 = io_read_0_addr[10] ? payload_10_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1639 = io_read_0_addr[11] ? payload_11_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1640 = io_read_0_addr[12] ? payload_12_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1641 = io_read_0_addr[13] ? payload_13_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1642 = io_read_0_addr[14] ? payload_14_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1643 = io_read_0_addr[15] ? payload_15_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1644 = _io_read_0_data_T_1628 | _io_read_0_data_T_1629; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1645 = _io_read_0_data_T_1644 | _io_read_0_data_T_1630; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1646 = _io_read_0_data_T_1645 | _io_read_0_data_T_1631; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1647 = _io_read_0_data_T_1646 | _io_read_0_data_T_1632; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1648 = _io_read_0_data_T_1647 | _io_read_0_data_T_1633; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1649 = _io_read_0_data_T_1648 | _io_read_0_data_T_1634; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1650 = _io_read_0_data_T_1649 | _io_read_0_data_T_1635; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1651 = _io_read_0_data_T_1650 | _io_read_0_data_T_1636; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1652 = _io_read_0_data_T_1651 | _io_read_0_data_T_1637; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1653 = _io_read_0_data_T_1652 | _io_read_0_data_T_1638; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1654 = _io_read_0_data_T_1653 | _io_read_0_data_T_1639; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1655 = _io_read_0_data_T_1654 | _io_read_0_data_T_1640; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1656 = _io_read_0_data_T_1655 | _io_read_0_data_T_1641; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_1657 = _io_read_0_data_T_1656 | _io_read_0_data_T_1642; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1907 = io_read_0_addr[0] ? payload_0_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1908 = io_read_0_addr[1] ? payload_1_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1909 = io_read_0_addr[2] ? payload_2_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1910 = io_read_0_addr[3] ? payload_3_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1911 = io_read_0_addr[4] ? payload_4_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1912 = io_read_0_addr[5] ? payload_5_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1913 = io_read_0_addr[6] ? payload_6_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1914 = io_read_0_addr[7] ? payload_7_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1915 = io_read_0_addr[8] ? payload_8_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1916 = io_read_0_addr[9] ? payload_9_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1917 = io_read_0_addr[10] ? payload_10_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1918 = io_read_0_addr[11] ? payload_11_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1919 = io_read_0_addr[12] ? payload_12_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1920 = io_read_0_addr[13] ? payload_13_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1921 = io_read_0_addr[14] ? payload_14_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1922 = io_read_0_addr[15] ? payload_15_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1923 = _io_read_0_data_T_1907 | _io_read_0_data_T_1908; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1924 = _io_read_0_data_T_1923 | _io_read_0_data_T_1909; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1925 = _io_read_0_data_T_1924 | _io_read_0_data_T_1910; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1926 = _io_read_0_data_T_1925 | _io_read_0_data_T_1911; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1927 = _io_read_0_data_T_1926 | _io_read_0_data_T_1912; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1928 = _io_read_0_data_T_1927 | _io_read_0_data_T_1913; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1929 = _io_read_0_data_T_1928 | _io_read_0_data_T_1914; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1930 = _io_read_0_data_T_1929 | _io_read_0_data_T_1915; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1931 = _io_read_0_data_T_1930 | _io_read_0_data_T_1916; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1932 = _io_read_0_data_T_1931 | _io_read_0_data_T_1917; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1933 = _io_read_0_data_T_1932 | _io_read_0_data_T_1918; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1934 = _io_read_0_data_T_1933 | _io_read_0_data_T_1919; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1935 = _io_read_0_data_T_1934 | _io_read_0_data_T_1920; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1936 = _io_read_0_data_T_1935 | _io_read_0_data_T_1921; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1938 = io_read_0_addr[0] ? payload_0_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1939 = io_read_0_addr[1] ? payload_1_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1940 = io_read_0_addr[2] ? payload_2_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1941 = io_read_0_addr[3] ? payload_3_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1942 = io_read_0_addr[4] ? payload_4_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1943 = io_read_0_addr[5] ? payload_5_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1944 = io_read_0_addr[6] ? payload_6_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1945 = io_read_0_addr[7] ? payload_7_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1946 = io_read_0_addr[8] ? payload_8_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1947 = io_read_0_addr[9] ? payload_9_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1948 = io_read_0_addr[10] ? payload_10_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1949 = io_read_0_addr[11] ? payload_11_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1950 = io_read_0_addr[12] ? payload_12_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1951 = io_read_0_addr[13] ? payload_13_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1952 = io_read_0_addr[14] ? payload_14_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1953 = io_read_0_addr[15] ? payload_15_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1954 = _io_read_0_data_T_1938 | _io_read_0_data_T_1939; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1955 = _io_read_0_data_T_1954 | _io_read_0_data_T_1940; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1956 = _io_read_0_data_T_1955 | _io_read_0_data_T_1941; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1957 = _io_read_0_data_T_1956 | _io_read_0_data_T_1942; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1958 = _io_read_0_data_T_1957 | _io_read_0_data_T_1943; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1959 = _io_read_0_data_T_1958 | _io_read_0_data_T_1944; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1960 = _io_read_0_data_T_1959 | _io_read_0_data_T_1945; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1961 = _io_read_0_data_T_1960 | _io_read_0_data_T_1946; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1962 = _io_read_0_data_T_1961 | _io_read_0_data_T_1947; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1963 = _io_read_0_data_T_1962 | _io_read_0_data_T_1948; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1964 = _io_read_0_data_T_1963 | _io_read_0_data_T_1949; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1965 = _io_read_0_data_T_1964 | _io_read_0_data_T_1950; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1966 = _io_read_0_data_T_1965 | _io_read_0_data_T_1951; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_1967 = _io_read_0_data_T_1966 | _io_read_0_data_T_1952; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_1984 = io_read_0_addr[15] & payload_15_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2000 = io_read_0_addr[0] ? payload_0_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2001 = io_read_0_addr[1] ? payload_1_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2002 = io_read_0_addr[2] ? payload_2_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2003 = io_read_0_addr[3] ? payload_3_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2004 = io_read_0_addr[4] ? payload_4_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2005 = io_read_0_addr[5] ? payload_5_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2006 = io_read_0_addr[6] ? payload_6_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2007 = io_read_0_addr[7] ? payload_7_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2008 = io_read_0_addr[8] ? payload_8_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2009 = io_read_0_addr[9] ? payload_9_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2010 = io_read_0_addr[10] ? payload_10_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2011 = io_read_0_addr[11] ? payload_11_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2012 = io_read_0_addr[12] ? payload_12_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2013 = io_read_0_addr[13] ? payload_13_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2014 = io_read_0_addr[14] ? payload_14_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2015 = io_read_0_addr[15] ? payload_15_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2016 = _io_read_0_data_T_2000 | _io_read_0_data_T_2001; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2017 = _io_read_0_data_T_2016 | _io_read_0_data_T_2002; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2018 = _io_read_0_data_T_2017 | _io_read_0_data_T_2003; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2019 = _io_read_0_data_T_2018 | _io_read_0_data_T_2004; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2020 = _io_read_0_data_T_2019 | _io_read_0_data_T_2005; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2021 = _io_read_0_data_T_2020 | _io_read_0_data_T_2006; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2022 = _io_read_0_data_T_2021 | _io_read_0_data_T_2007; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2023 = _io_read_0_data_T_2022 | _io_read_0_data_T_2008; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2024 = _io_read_0_data_T_2023 | _io_read_0_data_T_2009; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2025 = _io_read_0_data_T_2024 | _io_read_0_data_T_2010; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2026 = _io_read_0_data_T_2025 | _io_read_0_data_T_2011; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2027 = _io_read_0_data_T_2026 | _io_read_0_data_T_2012; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2028 = _io_read_0_data_T_2027 | _io_read_0_data_T_2013; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2029 = _io_read_0_data_T_2028 | _io_read_0_data_T_2014; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2046 = io_read_0_addr[15] & payload_15_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2077 = io_read_0_addr[15] & payload_15_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2093 = io_read_0_addr[0] ? payload_0_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2094 = io_read_0_addr[1] ? payload_1_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2095 = io_read_0_addr[2] ? payload_2_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2096 = io_read_0_addr[3] ? payload_3_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2097 = io_read_0_addr[4] ? payload_4_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2098 = io_read_0_addr[5] ? payload_5_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2099 = io_read_0_addr[6] ? payload_6_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2100 = io_read_0_addr[7] ? payload_7_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2101 = io_read_0_addr[8] ? payload_8_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2102 = io_read_0_addr[9] ? payload_9_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2103 = io_read_0_addr[10] ? payload_10_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2104 = io_read_0_addr[11] ? payload_11_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2105 = io_read_0_addr[12] ? payload_12_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2106 = io_read_0_addr[13] ? payload_13_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2107 = io_read_0_addr[14] ? payload_14_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2108 = io_read_0_addr[15] ? payload_15_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2109 = _io_read_0_data_T_2093 | _io_read_0_data_T_2094; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2110 = _io_read_0_data_T_2109 | _io_read_0_data_T_2095; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2111 = _io_read_0_data_T_2110 | _io_read_0_data_T_2096; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2112 = _io_read_0_data_T_2111 | _io_read_0_data_T_2097; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2113 = _io_read_0_data_T_2112 | _io_read_0_data_T_2098; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2114 = _io_read_0_data_T_2113 | _io_read_0_data_T_2099; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2115 = _io_read_0_data_T_2114 | _io_read_0_data_T_2100; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2116 = _io_read_0_data_T_2115 | _io_read_0_data_T_2101; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2117 = _io_read_0_data_T_2116 | _io_read_0_data_T_2102; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2118 = _io_read_0_data_T_2117 | _io_read_0_data_T_2103; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2119 = _io_read_0_data_T_2118 | _io_read_0_data_T_2104; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2120 = _io_read_0_data_T_2119 | _io_read_0_data_T_2105; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2121 = _io_read_0_data_T_2120 | _io_read_0_data_T_2106; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_2122 = _io_read_0_data_T_2121 | _io_read_0_data_T_2107; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2139 = io_read_0_addr[15] & payload_15_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2170 = io_read_0_addr[15] & payload_15_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2232 = io_read_0_addr[15] & payload_15_cf_pred_taken; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2263 = io_read_0_addr[15] & payload_15_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2294 = io_read_0_addr[15] & payload_15_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2310 = io_read_0_addr[0] ? payload_0_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2311 = io_read_0_addr[1] ? payload_1_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2312 = io_read_0_addr[2] ? payload_2_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2313 = io_read_0_addr[3] ? payload_3_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2314 = io_read_0_addr[4] ? payload_4_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2315 = io_read_0_addr[5] ? payload_5_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2316 = io_read_0_addr[6] ? payload_6_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2317 = io_read_0_addr[7] ? payload_7_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2318 = io_read_0_addr[8] ? payload_8_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2319 = io_read_0_addr[9] ? payload_9_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2320 = io_read_0_addr[10] ? payload_10_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2321 = io_read_0_addr[11] ? payload_11_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2322 = io_read_0_addr[12] ? payload_12_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2323 = io_read_0_addr[13] ? payload_13_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2324 = io_read_0_addr[14] ? payload_14_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2325 = io_read_0_addr[15] ? payload_15_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2326 = _io_read_0_data_T_2310 | _io_read_0_data_T_2311; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2327 = _io_read_0_data_T_2326 | _io_read_0_data_T_2312; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2328 = _io_read_0_data_T_2327 | _io_read_0_data_T_2313; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2329 = _io_read_0_data_T_2328 | _io_read_0_data_T_2314; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2330 = _io_read_0_data_T_2329 | _io_read_0_data_T_2315; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2331 = _io_read_0_data_T_2330 | _io_read_0_data_T_2316; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2332 = _io_read_0_data_T_2331 | _io_read_0_data_T_2317; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2333 = _io_read_0_data_T_2332 | _io_read_0_data_T_2318; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2334 = _io_read_0_data_T_2333 | _io_read_0_data_T_2319; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2335 = _io_read_0_data_T_2334 | _io_read_0_data_T_2320; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2336 = _io_read_0_data_T_2335 | _io_read_0_data_T_2321; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2337 = _io_read_0_data_T_2336 | _io_read_0_data_T_2322; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2338 = _io_read_0_data_T_2337 | _io_read_0_data_T_2323; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_2339 = _io_read_0_data_T_2338 | _io_read_0_data_T_2324; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2356 = io_read_0_addr[15] & payload_15_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2604 = io_read_0_addr[15] & payload_15_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  _io_read_0_data_T_2635 = io_read_0_addr[15] & payload_15_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3271 = io_read_0_addr[0] ? payload_0_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3272 = io_read_0_addr[1] ? payload_1_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3273 = io_read_0_addr[2] ? payload_2_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3274 = io_read_0_addr[3] ? payload_3_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3275 = io_read_0_addr[4] ? payload_4_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3276 = io_read_0_addr[5] ? payload_5_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3277 = io_read_0_addr[6] ? payload_6_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3278 = io_read_0_addr[7] ? payload_7_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3279 = io_read_0_addr[8] ? payload_8_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3280 = io_read_0_addr[9] ? payload_9_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3281 = io_read_0_addr[10] ? payload_10_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3282 = io_read_0_addr[11] ? payload_11_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3283 = io_read_0_addr[12] ? payload_12_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3284 = io_read_0_addr[13] ? payload_13_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3285 = io_read_0_addr[14] ? payload_14_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3286 = io_read_0_addr[15] ? payload_15_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3287 = _io_read_0_data_T_3271 | _io_read_0_data_T_3272; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3288 = _io_read_0_data_T_3287 | _io_read_0_data_T_3273; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3289 = _io_read_0_data_T_3288 | _io_read_0_data_T_3274; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3290 = _io_read_0_data_T_3289 | _io_read_0_data_T_3275; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3291 = _io_read_0_data_T_3290 | _io_read_0_data_T_3276; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3292 = _io_read_0_data_T_3291 | _io_read_0_data_T_3277; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3293 = _io_read_0_data_T_3292 | _io_read_0_data_T_3278; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3294 = _io_read_0_data_T_3293 | _io_read_0_data_T_3279; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3295 = _io_read_0_data_T_3294 | _io_read_0_data_T_3280; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3296 = _io_read_0_data_T_3295 | _io_read_0_data_T_3281; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3297 = _io_read_0_data_T_3296 | _io_read_0_data_T_3282; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3298 = _io_read_0_data_T_3297 | _io_read_0_data_T_3283; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3299 = _io_read_0_data_T_3298 | _io_read_0_data_T_3284; // @[Mux.scala 27:73]
  wire [9:0] _io_read_0_data_T_3300 = _io_read_0_data_T_3299 | _io_read_0_data_T_3285; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_357 = io_read_1_addr[0] ? payload_0_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_358 = io_read_1_addr[1] ? payload_1_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_359 = io_read_1_addr[2] ? payload_2_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_360 = io_read_1_addr[3] ? payload_3_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_361 = io_read_1_addr[4] ? payload_4_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_362 = io_read_1_addr[5] ? payload_5_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_363 = io_read_1_addr[6] ? payload_6_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_364 = io_read_1_addr[7] ? payload_7_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_365 = io_read_1_addr[8] ? payload_8_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_366 = io_read_1_addr[9] ? payload_9_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_367 = io_read_1_addr[10] ? payload_10_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_368 = io_read_1_addr[11] ? payload_11_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_369 = io_read_1_addr[12] ? payload_12_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_370 = io_read_1_addr[13] ? payload_13_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_371 = io_read_1_addr[14] ? payload_14_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_372 = io_read_1_addr[15] ? payload_15_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_373 = _io_read_1_data_T_357 | _io_read_1_data_T_358; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_374 = _io_read_1_data_T_373 | _io_read_1_data_T_359; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_375 = _io_read_1_data_T_374 | _io_read_1_data_T_360; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_376 = _io_read_1_data_T_375 | _io_read_1_data_T_361; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_377 = _io_read_1_data_T_376 | _io_read_1_data_T_362; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_378 = _io_read_1_data_T_377 | _io_read_1_data_T_363; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_379 = _io_read_1_data_T_378 | _io_read_1_data_T_364; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_380 = _io_read_1_data_T_379 | _io_read_1_data_T_365; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_381 = _io_read_1_data_T_380 | _io_read_1_data_T_366; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_382 = _io_read_1_data_T_381 | _io_read_1_data_T_367; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_383 = _io_read_1_data_T_382 | _io_read_1_data_T_368; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_384 = _io_read_1_data_T_383 | _io_read_1_data_T_369; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_385 = _io_read_1_data_T_384 | _io_read_1_data_T_370; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_386 = _io_read_1_data_T_385 | _io_read_1_data_T_371; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_403 = io_read_1_addr[15] & payload_15_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_419 = io_read_1_addr[0] ? payload_0_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_420 = io_read_1_addr[1] ? payload_1_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_421 = io_read_1_addr[2] ? payload_2_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_422 = io_read_1_addr[3] ? payload_3_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_423 = io_read_1_addr[4] ? payload_4_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_424 = io_read_1_addr[5] ? payload_5_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_425 = io_read_1_addr[6] ? payload_6_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_426 = io_read_1_addr[7] ? payload_7_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_427 = io_read_1_addr[8] ? payload_8_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_428 = io_read_1_addr[9] ? payload_9_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_429 = io_read_1_addr[10] ? payload_10_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_430 = io_read_1_addr[11] ? payload_11_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_431 = io_read_1_addr[12] ? payload_12_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_432 = io_read_1_addr[13] ? payload_13_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_433 = io_read_1_addr[14] ? payload_14_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_434 = io_read_1_addr[15] ? payload_15_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_435 = _io_read_1_data_T_419 | _io_read_1_data_T_420; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_436 = _io_read_1_data_T_435 | _io_read_1_data_T_421; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_437 = _io_read_1_data_T_436 | _io_read_1_data_T_422; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_438 = _io_read_1_data_T_437 | _io_read_1_data_T_423; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_439 = _io_read_1_data_T_438 | _io_read_1_data_T_424; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_440 = _io_read_1_data_T_439 | _io_read_1_data_T_425; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_441 = _io_read_1_data_T_440 | _io_read_1_data_T_426; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_442 = _io_read_1_data_T_441 | _io_read_1_data_T_427; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_443 = _io_read_1_data_T_442 | _io_read_1_data_T_428; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_444 = _io_read_1_data_T_443 | _io_read_1_data_T_429; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_445 = _io_read_1_data_T_444 | _io_read_1_data_T_430; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_446 = _io_read_1_data_T_445 | _io_read_1_data_T_431; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_447 = _io_read_1_data_T_446 | _io_read_1_data_T_432; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_448 = _io_read_1_data_T_447 | _io_read_1_data_T_433; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_465 = io_read_1_addr[15] & payload_15_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_481 = io_read_1_addr[0] ? payload_0_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_482 = io_read_1_addr[1] ? payload_1_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_483 = io_read_1_addr[2] ? payload_2_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_484 = io_read_1_addr[3] ? payload_3_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_485 = io_read_1_addr[4] ? payload_4_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_486 = io_read_1_addr[5] ? payload_5_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_487 = io_read_1_addr[6] ? payload_6_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_488 = io_read_1_addr[7] ? payload_7_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_489 = io_read_1_addr[8] ? payload_8_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_490 = io_read_1_addr[9] ? payload_9_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_491 = io_read_1_addr[10] ? payload_10_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_492 = io_read_1_addr[11] ? payload_11_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_493 = io_read_1_addr[12] ? payload_12_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_494 = io_read_1_addr[13] ? payload_13_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_495 = io_read_1_addr[14] ? payload_14_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_496 = io_read_1_addr[15] ? payload_15_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_497 = _io_read_1_data_T_481 | _io_read_1_data_T_482; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_498 = _io_read_1_data_T_497 | _io_read_1_data_T_483; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_499 = _io_read_1_data_T_498 | _io_read_1_data_T_484; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_500 = _io_read_1_data_T_499 | _io_read_1_data_T_485; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_501 = _io_read_1_data_T_500 | _io_read_1_data_T_486; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_502 = _io_read_1_data_T_501 | _io_read_1_data_T_487; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_503 = _io_read_1_data_T_502 | _io_read_1_data_T_488; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_504 = _io_read_1_data_T_503 | _io_read_1_data_T_489; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_505 = _io_read_1_data_T_504 | _io_read_1_data_T_490; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_506 = _io_read_1_data_T_505 | _io_read_1_data_T_491; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_507 = _io_read_1_data_T_506 | _io_read_1_data_T_492; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_508 = _io_read_1_data_T_507 | _io_read_1_data_T_493; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_509 = _io_read_1_data_T_508 | _io_read_1_data_T_494; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_510 = _io_read_1_data_T_509 | _io_read_1_data_T_495; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_527 = io_read_1_addr[15] & payload_15_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_574 = io_read_1_addr[0] ? payload_0_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_575 = io_read_1_addr[1] ? payload_1_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_576 = io_read_1_addr[2] ? payload_2_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_577 = io_read_1_addr[3] ? payload_3_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_578 = io_read_1_addr[4] ? payload_4_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_579 = io_read_1_addr[5] ? payload_5_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_580 = io_read_1_addr[6] ? payload_6_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_581 = io_read_1_addr[7] ? payload_7_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_582 = io_read_1_addr[8] ? payload_8_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_583 = io_read_1_addr[9] ? payload_9_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_584 = io_read_1_addr[10] ? payload_10_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_585 = io_read_1_addr[11] ? payload_11_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_586 = io_read_1_addr[12] ? payload_12_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_587 = io_read_1_addr[13] ? payload_13_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_588 = io_read_1_addr[14] ? payload_14_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_589 = io_read_1_addr[15] ? payload_15_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_590 = _io_read_1_data_T_574 | _io_read_1_data_T_575; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_591 = _io_read_1_data_T_590 | _io_read_1_data_T_576; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_592 = _io_read_1_data_T_591 | _io_read_1_data_T_577; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_593 = _io_read_1_data_T_592 | _io_read_1_data_T_578; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_594 = _io_read_1_data_T_593 | _io_read_1_data_T_579; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_595 = _io_read_1_data_T_594 | _io_read_1_data_T_580; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_596 = _io_read_1_data_T_595 | _io_read_1_data_T_581; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_597 = _io_read_1_data_T_596 | _io_read_1_data_T_582; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_598 = _io_read_1_data_T_597 | _io_read_1_data_T_583; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_599 = _io_read_1_data_T_598 | _io_read_1_data_T_584; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_600 = _io_read_1_data_T_599 | _io_read_1_data_T_585; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_601 = _io_read_1_data_T_600 | _io_read_1_data_T_586; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_602 = _io_read_1_data_T_601 | _io_read_1_data_T_587; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_603 = _io_read_1_data_T_602 | _io_read_1_data_T_588; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1349 = io_read_1_addr[0] ? payload_0_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1350 = io_read_1_addr[1] ? payload_1_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1351 = io_read_1_addr[2] ? payload_2_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1352 = io_read_1_addr[3] ? payload_3_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1353 = io_read_1_addr[4] ? payload_4_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1354 = io_read_1_addr[5] ? payload_5_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1355 = io_read_1_addr[6] ? payload_6_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1356 = io_read_1_addr[7] ? payload_7_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1357 = io_read_1_addr[8] ? payload_8_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1358 = io_read_1_addr[9] ? payload_9_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1359 = io_read_1_addr[10] ? payload_10_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1360 = io_read_1_addr[11] ? payload_11_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1361 = io_read_1_addr[12] ? payload_12_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1362 = io_read_1_addr[13] ? payload_13_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1363 = io_read_1_addr[14] ? payload_14_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1364 = io_read_1_addr[15] ? payload_15_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1365 = _io_read_1_data_T_1349 | _io_read_1_data_T_1350; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1366 = _io_read_1_data_T_1365 | _io_read_1_data_T_1351; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1367 = _io_read_1_data_T_1366 | _io_read_1_data_T_1352; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1368 = _io_read_1_data_T_1367 | _io_read_1_data_T_1353; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1369 = _io_read_1_data_T_1368 | _io_read_1_data_T_1354; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1370 = _io_read_1_data_T_1369 | _io_read_1_data_T_1355; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1371 = _io_read_1_data_T_1370 | _io_read_1_data_T_1356; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1372 = _io_read_1_data_T_1371 | _io_read_1_data_T_1357; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1373 = _io_read_1_data_T_1372 | _io_read_1_data_T_1358; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1374 = _io_read_1_data_T_1373 | _io_read_1_data_T_1359; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1375 = _io_read_1_data_T_1374 | _io_read_1_data_T_1360; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1376 = _io_read_1_data_T_1375 | _io_read_1_data_T_1361; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1377 = _io_read_1_data_T_1376 | _io_read_1_data_T_1362; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_1378 = _io_read_1_data_T_1377 | _io_read_1_data_T_1363; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_1550 = io_read_1_addr[15] & payload_15_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_1581 = io_read_1_addr[15] & payload_15_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1597 = io_read_1_addr[0] ? payload_0_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1598 = io_read_1_addr[1] ? payload_1_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1599 = io_read_1_addr[2] ? payload_2_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1600 = io_read_1_addr[3] ? payload_3_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1601 = io_read_1_addr[4] ? payload_4_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1602 = io_read_1_addr[5] ? payload_5_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1603 = io_read_1_addr[6] ? payload_6_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1604 = io_read_1_addr[7] ? payload_7_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1605 = io_read_1_addr[8] ? payload_8_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1606 = io_read_1_addr[9] ? payload_9_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1607 = io_read_1_addr[10] ? payload_10_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1608 = io_read_1_addr[11] ? payload_11_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1609 = io_read_1_addr[12] ? payload_12_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1610 = io_read_1_addr[13] ? payload_13_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1611 = io_read_1_addr[14] ? payload_14_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1612 = io_read_1_addr[15] ? payload_15_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1613 = _io_read_1_data_T_1597 | _io_read_1_data_T_1598; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1614 = _io_read_1_data_T_1613 | _io_read_1_data_T_1599; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1615 = _io_read_1_data_T_1614 | _io_read_1_data_T_1600; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1616 = _io_read_1_data_T_1615 | _io_read_1_data_T_1601; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1617 = _io_read_1_data_T_1616 | _io_read_1_data_T_1602; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1618 = _io_read_1_data_T_1617 | _io_read_1_data_T_1603; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1619 = _io_read_1_data_T_1618 | _io_read_1_data_T_1604; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1620 = _io_read_1_data_T_1619 | _io_read_1_data_T_1605; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1621 = _io_read_1_data_T_1620 | _io_read_1_data_T_1606; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1622 = _io_read_1_data_T_1621 | _io_read_1_data_T_1607; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1623 = _io_read_1_data_T_1622 | _io_read_1_data_T_1608; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1624 = _io_read_1_data_T_1623 | _io_read_1_data_T_1609; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1625 = _io_read_1_data_T_1624 | _io_read_1_data_T_1610; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_1626 = _io_read_1_data_T_1625 | _io_read_1_data_T_1611; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1628 = io_read_1_addr[0] ? payload_0_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1629 = io_read_1_addr[1] ? payload_1_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1630 = io_read_1_addr[2] ? payload_2_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1631 = io_read_1_addr[3] ? payload_3_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1632 = io_read_1_addr[4] ? payload_4_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1633 = io_read_1_addr[5] ? payload_5_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1634 = io_read_1_addr[6] ? payload_6_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1635 = io_read_1_addr[7] ? payload_7_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1636 = io_read_1_addr[8] ? payload_8_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1637 = io_read_1_addr[9] ? payload_9_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1638 = io_read_1_addr[10] ? payload_10_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1639 = io_read_1_addr[11] ? payload_11_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1640 = io_read_1_addr[12] ? payload_12_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1641 = io_read_1_addr[13] ? payload_13_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1642 = io_read_1_addr[14] ? payload_14_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1643 = io_read_1_addr[15] ? payload_15_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1644 = _io_read_1_data_T_1628 | _io_read_1_data_T_1629; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1645 = _io_read_1_data_T_1644 | _io_read_1_data_T_1630; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1646 = _io_read_1_data_T_1645 | _io_read_1_data_T_1631; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1647 = _io_read_1_data_T_1646 | _io_read_1_data_T_1632; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1648 = _io_read_1_data_T_1647 | _io_read_1_data_T_1633; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1649 = _io_read_1_data_T_1648 | _io_read_1_data_T_1634; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1650 = _io_read_1_data_T_1649 | _io_read_1_data_T_1635; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1651 = _io_read_1_data_T_1650 | _io_read_1_data_T_1636; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1652 = _io_read_1_data_T_1651 | _io_read_1_data_T_1637; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1653 = _io_read_1_data_T_1652 | _io_read_1_data_T_1638; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1654 = _io_read_1_data_T_1653 | _io_read_1_data_T_1639; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1655 = _io_read_1_data_T_1654 | _io_read_1_data_T_1640; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1656 = _io_read_1_data_T_1655 | _io_read_1_data_T_1641; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_1657 = _io_read_1_data_T_1656 | _io_read_1_data_T_1642; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1907 = io_read_1_addr[0] ? payload_0_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1908 = io_read_1_addr[1] ? payload_1_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1909 = io_read_1_addr[2] ? payload_2_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1910 = io_read_1_addr[3] ? payload_3_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1911 = io_read_1_addr[4] ? payload_4_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1912 = io_read_1_addr[5] ? payload_5_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1913 = io_read_1_addr[6] ? payload_6_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1914 = io_read_1_addr[7] ? payload_7_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1915 = io_read_1_addr[8] ? payload_8_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1916 = io_read_1_addr[9] ? payload_9_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1917 = io_read_1_addr[10] ? payload_10_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1918 = io_read_1_addr[11] ? payload_11_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1919 = io_read_1_addr[12] ? payload_12_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1920 = io_read_1_addr[13] ? payload_13_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1921 = io_read_1_addr[14] ? payload_14_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1922 = io_read_1_addr[15] ? payload_15_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1923 = _io_read_1_data_T_1907 | _io_read_1_data_T_1908; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1924 = _io_read_1_data_T_1923 | _io_read_1_data_T_1909; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1925 = _io_read_1_data_T_1924 | _io_read_1_data_T_1910; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1926 = _io_read_1_data_T_1925 | _io_read_1_data_T_1911; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1927 = _io_read_1_data_T_1926 | _io_read_1_data_T_1912; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1928 = _io_read_1_data_T_1927 | _io_read_1_data_T_1913; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1929 = _io_read_1_data_T_1928 | _io_read_1_data_T_1914; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1930 = _io_read_1_data_T_1929 | _io_read_1_data_T_1915; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1931 = _io_read_1_data_T_1930 | _io_read_1_data_T_1916; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1932 = _io_read_1_data_T_1931 | _io_read_1_data_T_1917; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1933 = _io_read_1_data_T_1932 | _io_read_1_data_T_1918; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1934 = _io_read_1_data_T_1933 | _io_read_1_data_T_1919; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1935 = _io_read_1_data_T_1934 | _io_read_1_data_T_1920; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1936 = _io_read_1_data_T_1935 | _io_read_1_data_T_1921; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1938 = io_read_1_addr[0] ? payload_0_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1939 = io_read_1_addr[1] ? payload_1_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1940 = io_read_1_addr[2] ? payload_2_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1941 = io_read_1_addr[3] ? payload_3_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1942 = io_read_1_addr[4] ? payload_4_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1943 = io_read_1_addr[5] ? payload_5_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1944 = io_read_1_addr[6] ? payload_6_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1945 = io_read_1_addr[7] ? payload_7_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1946 = io_read_1_addr[8] ? payload_8_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1947 = io_read_1_addr[9] ? payload_9_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1948 = io_read_1_addr[10] ? payload_10_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1949 = io_read_1_addr[11] ? payload_11_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1950 = io_read_1_addr[12] ? payload_12_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1951 = io_read_1_addr[13] ? payload_13_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1952 = io_read_1_addr[14] ? payload_14_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1953 = io_read_1_addr[15] ? payload_15_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1954 = _io_read_1_data_T_1938 | _io_read_1_data_T_1939; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1955 = _io_read_1_data_T_1954 | _io_read_1_data_T_1940; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1956 = _io_read_1_data_T_1955 | _io_read_1_data_T_1941; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1957 = _io_read_1_data_T_1956 | _io_read_1_data_T_1942; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1958 = _io_read_1_data_T_1957 | _io_read_1_data_T_1943; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1959 = _io_read_1_data_T_1958 | _io_read_1_data_T_1944; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1960 = _io_read_1_data_T_1959 | _io_read_1_data_T_1945; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1961 = _io_read_1_data_T_1960 | _io_read_1_data_T_1946; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1962 = _io_read_1_data_T_1961 | _io_read_1_data_T_1947; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1963 = _io_read_1_data_T_1962 | _io_read_1_data_T_1948; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1964 = _io_read_1_data_T_1963 | _io_read_1_data_T_1949; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1965 = _io_read_1_data_T_1964 | _io_read_1_data_T_1950; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1966 = _io_read_1_data_T_1965 | _io_read_1_data_T_1951; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_1967 = _io_read_1_data_T_1966 | _io_read_1_data_T_1952; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_1984 = io_read_1_addr[15] & payload_15_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2000 = io_read_1_addr[0] ? payload_0_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2001 = io_read_1_addr[1] ? payload_1_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2002 = io_read_1_addr[2] ? payload_2_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2003 = io_read_1_addr[3] ? payload_3_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2004 = io_read_1_addr[4] ? payload_4_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2005 = io_read_1_addr[5] ? payload_5_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2006 = io_read_1_addr[6] ? payload_6_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2007 = io_read_1_addr[7] ? payload_7_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2008 = io_read_1_addr[8] ? payload_8_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2009 = io_read_1_addr[9] ? payload_9_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2010 = io_read_1_addr[10] ? payload_10_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2011 = io_read_1_addr[11] ? payload_11_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2012 = io_read_1_addr[12] ? payload_12_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2013 = io_read_1_addr[13] ? payload_13_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2014 = io_read_1_addr[14] ? payload_14_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2015 = io_read_1_addr[15] ? payload_15_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2016 = _io_read_1_data_T_2000 | _io_read_1_data_T_2001; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2017 = _io_read_1_data_T_2016 | _io_read_1_data_T_2002; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2018 = _io_read_1_data_T_2017 | _io_read_1_data_T_2003; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2019 = _io_read_1_data_T_2018 | _io_read_1_data_T_2004; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2020 = _io_read_1_data_T_2019 | _io_read_1_data_T_2005; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2021 = _io_read_1_data_T_2020 | _io_read_1_data_T_2006; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2022 = _io_read_1_data_T_2021 | _io_read_1_data_T_2007; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2023 = _io_read_1_data_T_2022 | _io_read_1_data_T_2008; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2024 = _io_read_1_data_T_2023 | _io_read_1_data_T_2009; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2025 = _io_read_1_data_T_2024 | _io_read_1_data_T_2010; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2026 = _io_read_1_data_T_2025 | _io_read_1_data_T_2011; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2027 = _io_read_1_data_T_2026 | _io_read_1_data_T_2012; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2028 = _io_read_1_data_T_2027 | _io_read_1_data_T_2013; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2029 = _io_read_1_data_T_2028 | _io_read_1_data_T_2014; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2046 = io_read_1_addr[15] & payload_15_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2077 = io_read_1_addr[15] & payload_15_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2093 = io_read_1_addr[0] ? payload_0_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2094 = io_read_1_addr[1] ? payload_1_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2095 = io_read_1_addr[2] ? payload_2_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2096 = io_read_1_addr[3] ? payload_3_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2097 = io_read_1_addr[4] ? payload_4_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2098 = io_read_1_addr[5] ? payload_5_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2099 = io_read_1_addr[6] ? payload_6_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2100 = io_read_1_addr[7] ? payload_7_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2101 = io_read_1_addr[8] ? payload_8_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2102 = io_read_1_addr[9] ? payload_9_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2103 = io_read_1_addr[10] ? payload_10_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2104 = io_read_1_addr[11] ? payload_11_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2105 = io_read_1_addr[12] ? payload_12_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2106 = io_read_1_addr[13] ? payload_13_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2107 = io_read_1_addr[14] ? payload_14_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2108 = io_read_1_addr[15] ? payload_15_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2109 = _io_read_1_data_T_2093 | _io_read_1_data_T_2094; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2110 = _io_read_1_data_T_2109 | _io_read_1_data_T_2095; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2111 = _io_read_1_data_T_2110 | _io_read_1_data_T_2096; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2112 = _io_read_1_data_T_2111 | _io_read_1_data_T_2097; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2113 = _io_read_1_data_T_2112 | _io_read_1_data_T_2098; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2114 = _io_read_1_data_T_2113 | _io_read_1_data_T_2099; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2115 = _io_read_1_data_T_2114 | _io_read_1_data_T_2100; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2116 = _io_read_1_data_T_2115 | _io_read_1_data_T_2101; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2117 = _io_read_1_data_T_2116 | _io_read_1_data_T_2102; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2118 = _io_read_1_data_T_2117 | _io_read_1_data_T_2103; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2119 = _io_read_1_data_T_2118 | _io_read_1_data_T_2104; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2120 = _io_read_1_data_T_2119 | _io_read_1_data_T_2105; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2121 = _io_read_1_data_T_2120 | _io_read_1_data_T_2106; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_2122 = _io_read_1_data_T_2121 | _io_read_1_data_T_2107; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2139 = io_read_1_addr[15] & payload_15_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2170 = io_read_1_addr[15] & payload_15_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2232 = io_read_1_addr[15] & payload_15_cf_pred_taken; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2263 = io_read_1_addr[15] & payload_15_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2294 = io_read_1_addr[15] & payload_15_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2310 = io_read_1_addr[0] ? payload_0_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2311 = io_read_1_addr[1] ? payload_1_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2312 = io_read_1_addr[2] ? payload_2_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2313 = io_read_1_addr[3] ? payload_3_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2314 = io_read_1_addr[4] ? payload_4_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2315 = io_read_1_addr[5] ? payload_5_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2316 = io_read_1_addr[6] ? payload_6_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2317 = io_read_1_addr[7] ? payload_7_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2318 = io_read_1_addr[8] ? payload_8_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2319 = io_read_1_addr[9] ? payload_9_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2320 = io_read_1_addr[10] ? payload_10_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2321 = io_read_1_addr[11] ? payload_11_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2322 = io_read_1_addr[12] ? payload_12_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2323 = io_read_1_addr[13] ? payload_13_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2324 = io_read_1_addr[14] ? payload_14_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2325 = io_read_1_addr[15] ? payload_15_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2326 = _io_read_1_data_T_2310 | _io_read_1_data_T_2311; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2327 = _io_read_1_data_T_2326 | _io_read_1_data_T_2312; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2328 = _io_read_1_data_T_2327 | _io_read_1_data_T_2313; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2329 = _io_read_1_data_T_2328 | _io_read_1_data_T_2314; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2330 = _io_read_1_data_T_2329 | _io_read_1_data_T_2315; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2331 = _io_read_1_data_T_2330 | _io_read_1_data_T_2316; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2332 = _io_read_1_data_T_2331 | _io_read_1_data_T_2317; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2333 = _io_read_1_data_T_2332 | _io_read_1_data_T_2318; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2334 = _io_read_1_data_T_2333 | _io_read_1_data_T_2319; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2335 = _io_read_1_data_T_2334 | _io_read_1_data_T_2320; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2336 = _io_read_1_data_T_2335 | _io_read_1_data_T_2321; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2337 = _io_read_1_data_T_2336 | _io_read_1_data_T_2322; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2338 = _io_read_1_data_T_2337 | _io_read_1_data_T_2323; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_2339 = _io_read_1_data_T_2338 | _io_read_1_data_T_2324; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2356 = io_read_1_addr[15] & payload_15_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2604 = io_read_1_addr[15] & payload_15_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  _io_read_1_data_T_2635 = io_read_1_addr[15] & payload_15_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3271 = io_read_1_addr[0] ? payload_0_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3272 = io_read_1_addr[1] ? payload_1_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3273 = io_read_1_addr[2] ? payload_2_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3274 = io_read_1_addr[3] ? payload_3_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3275 = io_read_1_addr[4] ? payload_4_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3276 = io_read_1_addr[5] ? payload_5_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3277 = io_read_1_addr[6] ? payload_6_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3278 = io_read_1_addr[7] ? payload_7_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3279 = io_read_1_addr[8] ? payload_8_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3280 = io_read_1_addr[9] ? payload_9_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3281 = io_read_1_addr[10] ? payload_10_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3282 = io_read_1_addr[11] ? payload_11_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3283 = io_read_1_addr[12] ? payload_12_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3284 = io_read_1_addr[13] ? payload_13_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3285 = io_read_1_addr[14] ? payload_14_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3286 = io_read_1_addr[15] ? payload_15_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3287 = _io_read_1_data_T_3271 | _io_read_1_data_T_3272; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3288 = _io_read_1_data_T_3287 | _io_read_1_data_T_3273; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3289 = _io_read_1_data_T_3288 | _io_read_1_data_T_3274; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3290 = _io_read_1_data_T_3289 | _io_read_1_data_T_3275; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3291 = _io_read_1_data_T_3290 | _io_read_1_data_T_3276; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3292 = _io_read_1_data_T_3291 | _io_read_1_data_T_3277; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3293 = _io_read_1_data_T_3292 | _io_read_1_data_T_3278; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3294 = _io_read_1_data_T_3293 | _io_read_1_data_T_3279; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3295 = _io_read_1_data_T_3294 | _io_read_1_data_T_3280; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3296 = _io_read_1_data_T_3295 | _io_read_1_data_T_3281; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3297 = _io_read_1_data_T_3296 | _io_read_1_data_T_3282; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3298 = _io_read_1_data_T_3297 | _io_read_1_data_T_3283; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3299 = _io_read_1_data_T_3298 | _io_read_1_data_T_3284; // @[Mux.scala 27:73]
  wire [9:0] _io_read_1_data_T_3300 = _io_read_1_data_T_3299 | _io_read_1_data_T_3285; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_357 = io_read_2_addr[0] ? payload_0_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_358 = io_read_2_addr[1] ? payload_1_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_359 = io_read_2_addr[2] ? payload_2_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_360 = io_read_2_addr[3] ? payload_3_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_361 = io_read_2_addr[4] ? payload_4_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_362 = io_read_2_addr[5] ? payload_5_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_363 = io_read_2_addr[6] ? payload_6_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_364 = io_read_2_addr[7] ? payload_7_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_365 = io_read_2_addr[8] ? payload_8_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_366 = io_read_2_addr[9] ? payload_9_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_367 = io_read_2_addr[10] ? payload_10_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_368 = io_read_2_addr[11] ? payload_11_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_369 = io_read_2_addr[12] ? payload_12_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_370 = io_read_2_addr[13] ? payload_13_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_371 = io_read_2_addr[14] ? payload_14_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_372 = io_read_2_addr[15] ? payload_15_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_373 = _io_read_2_data_T_357 | _io_read_2_data_T_358; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_374 = _io_read_2_data_T_373 | _io_read_2_data_T_359; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_375 = _io_read_2_data_T_374 | _io_read_2_data_T_360; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_376 = _io_read_2_data_T_375 | _io_read_2_data_T_361; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_377 = _io_read_2_data_T_376 | _io_read_2_data_T_362; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_378 = _io_read_2_data_T_377 | _io_read_2_data_T_363; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_379 = _io_read_2_data_T_378 | _io_read_2_data_T_364; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_380 = _io_read_2_data_T_379 | _io_read_2_data_T_365; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_381 = _io_read_2_data_T_380 | _io_read_2_data_T_366; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_382 = _io_read_2_data_T_381 | _io_read_2_data_T_367; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_383 = _io_read_2_data_T_382 | _io_read_2_data_T_368; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_384 = _io_read_2_data_T_383 | _io_read_2_data_T_369; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_385 = _io_read_2_data_T_384 | _io_read_2_data_T_370; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_386 = _io_read_2_data_T_385 | _io_read_2_data_T_371; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_403 = io_read_2_addr[15] & payload_15_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_419 = io_read_2_addr[0] ? payload_0_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_420 = io_read_2_addr[1] ? payload_1_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_421 = io_read_2_addr[2] ? payload_2_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_422 = io_read_2_addr[3] ? payload_3_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_423 = io_read_2_addr[4] ? payload_4_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_424 = io_read_2_addr[5] ? payload_5_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_425 = io_read_2_addr[6] ? payload_6_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_426 = io_read_2_addr[7] ? payload_7_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_427 = io_read_2_addr[8] ? payload_8_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_428 = io_read_2_addr[9] ? payload_9_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_429 = io_read_2_addr[10] ? payload_10_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_430 = io_read_2_addr[11] ? payload_11_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_431 = io_read_2_addr[12] ? payload_12_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_432 = io_read_2_addr[13] ? payload_13_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_433 = io_read_2_addr[14] ? payload_14_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_434 = io_read_2_addr[15] ? payload_15_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_435 = _io_read_2_data_T_419 | _io_read_2_data_T_420; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_436 = _io_read_2_data_T_435 | _io_read_2_data_T_421; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_437 = _io_read_2_data_T_436 | _io_read_2_data_T_422; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_438 = _io_read_2_data_T_437 | _io_read_2_data_T_423; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_439 = _io_read_2_data_T_438 | _io_read_2_data_T_424; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_440 = _io_read_2_data_T_439 | _io_read_2_data_T_425; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_441 = _io_read_2_data_T_440 | _io_read_2_data_T_426; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_442 = _io_read_2_data_T_441 | _io_read_2_data_T_427; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_443 = _io_read_2_data_T_442 | _io_read_2_data_T_428; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_444 = _io_read_2_data_T_443 | _io_read_2_data_T_429; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_445 = _io_read_2_data_T_444 | _io_read_2_data_T_430; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_446 = _io_read_2_data_T_445 | _io_read_2_data_T_431; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_447 = _io_read_2_data_T_446 | _io_read_2_data_T_432; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_448 = _io_read_2_data_T_447 | _io_read_2_data_T_433; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_465 = io_read_2_addr[15] & payload_15_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_481 = io_read_2_addr[0] ? payload_0_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_482 = io_read_2_addr[1] ? payload_1_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_483 = io_read_2_addr[2] ? payload_2_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_484 = io_read_2_addr[3] ? payload_3_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_485 = io_read_2_addr[4] ? payload_4_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_486 = io_read_2_addr[5] ? payload_5_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_487 = io_read_2_addr[6] ? payload_6_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_488 = io_read_2_addr[7] ? payload_7_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_489 = io_read_2_addr[8] ? payload_8_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_490 = io_read_2_addr[9] ? payload_9_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_491 = io_read_2_addr[10] ? payload_10_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_492 = io_read_2_addr[11] ? payload_11_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_493 = io_read_2_addr[12] ? payload_12_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_494 = io_read_2_addr[13] ? payload_13_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_495 = io_read_2_addr[14] ? payload_14_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_496 = io_read_2_addr[15] ? payload_15_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_497 = _io_read_2_data_T_481 | _io_read_2_data_T_482; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_498 = _io_read_2_data_T_497 | _io_read_2_data_T_483; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_499 = _io_read_2_data_T_498 | _io_read_2_data_T_484; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_500 = _io_read_2_data_T_499 | _io_read_2_data_T_485; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_501 = _io_read_2_data_T_500 | _io_read_2_data_T_486; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_502 = _io_read_2_data_T_501 | _io_read_2_data_T_487; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_503 = _io_read_2_data_T_502 | _io_read_2_data_T_488; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_504 = _io_read_2_data_T_503 | _io_read_2_data_T_489; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_505 = _io_read_2_data_T_504 | _io_read_2_data_T_490; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_506 = _io_read_2_data_T_505 | _io_read_2_data_T_491; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_507 = _io_read_2_data_T_506 | _io_read_2_data_T_492; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_508 = _io_read_2_data_T_507 | _io_read_2_data_T_493; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_509 = _io_read_2_data_T_508 | _io_read_2_data_T_494; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_510 = _io_read_2_data_T_509 | _io_read_2_data_T_495; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_527 = io_read_2_addr[15] & payload_15_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_574 = io_read_2_addr[0] ? payload_0_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_575 = io_read_2_addr[1] ? payload_1_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_576 = io_read_2_addr[2] ? payload_2_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_577 = io_read_2_addr[3] ? payload_3_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_578 = io_read_2_addr[4] ? payload_4_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_579 = io_read_2_addr[5] ? payload_5_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_580 = io_read_2_addr[6] ? payload_6_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_581 = io_read_2_addr[7] ? payload_7_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_582 = io_read_2_addr[8] ? payload_8_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_583 = io_read_2_addr[9] ? payload_9_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_584 = io_read_2_addr[10] ? payload_10_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_585 = io_read_2_addr[11] ? payload_11_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_586 = io_read_2_addr[12] ? payload_12_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_587 = io_read_2_addr[13] ? payload_13_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_588 = io_read_2_addr[14] ? payload_14_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_589 = io_read_2_addr[15] ? payload_15_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_590 = _io_read_2_data_T_574 | _io_read_2_data_T_575; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_591 = _io_read_2_data_T_590 | _io_read_2_data_T_576; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_592 = _io_read_2_data_T_591 | _io_read_2_data_T_577; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_593 = _io_read_2_data_T_592 | _io_read_2_data_T_578; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_594 = _io_read_2_data_T_593 | _io_read_2_data_T_579; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_595 = _io_read_2_data_T_594 | _io_read_2_data_T_580; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_596 = _io_read_2_data_T_595 | _io_read_2_data_T_581; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_597 = _io_read_2_data_T_596 | _io_read_2_data_T_582; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_598 = _io_read_2_data_T_597 | _io_read_2_data_T_583; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_599 = _io_read_2_data_T_598 | _io_read_2_data_T_584; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_600 = _io_read_2_data_T_599 | _io_read_2_data_T_585; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_601 = _io_read_2_data_T_600 | _io_read_2_data_T_586; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_602 = _io_read_2_data_T_601 | _io_read_2_data_T_587; // @[Mux.scala 27:73]
  wire [5:0] _io_read_2_data_T_603 = _io_read_2_data_T_602 | _io_read_2_data_T_588; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1349 = io_read_2_addr[0] ? payload_0_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1350 = io_read_2_addr[1] ? payload_1_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1351 = io_read_2_addr[2] ? payload_2_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1352 = io_read_2_addr[3] ? payload_3_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1353 = io_read_2_addr[4] ? payload_4_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1354 = io_read_2_addr[5] ? payload_5_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1355 = io_read_2_addr[6] ? payload_6_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1356 = io_read_2_addr[7] ? payload_7_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1357 = io_read_2_addr[8] ? payload_8_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1358 = io_read_2_addr[9] ? payload_9_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1359 = io_read_2_addr[10] ? payload_10_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1360 = io_read_2_addr[11] ? payload_11_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1361 = io_read_2_addr[12] ? payload_12_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1362 = io_read_2_addr[13] ? payload_13_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1363 = io_read_2_addr[14] ? payload_14_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1364 = io_read_2_addr[15] ? payload_15_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1365 = _io_read_2_data_T_1349 | _io_read_2_data_T_1350; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1366 = _io_read_2_data_T_1365 | _io_read_2_data_T_1351; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1367 = _io_read_2_data_T_1366 | _io_read_2_data_T_1352; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1368 = _io_read_2_data_T_1367 | _io_read_2_data_T_1353; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1369 = _io_read_2_data_T_1368 | _io_read_2_data_T_1354; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1370 = _io_read_2_data_T_1369 | _io_read_2_data_T_1355; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1371 = _io_read_2_data_T_1370 | _io_read_2_data_T_1356; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1372 = _io_read_2_data_T_1371 | _io_read_2_data_T_1357; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1373 = _io_read_2_data_T_1372 | _io_read_2_data_T_1358; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1374 = _io_read_2_data_T_1373 | _io_read_2_data_T_1359; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1375 = _io_read_2_data_T_1374 | _io_read_2_data_T_1360; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1376 = _io_read_2_data_T_1375 | _io_read_2_data_T_1361; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1377 = _io_read_2_data_T_1376 | _io_read_2_data_T_1362; // @[Mux.scala 27:73]
  wire [19:0] _io_read_2_data_T_1378 = _io_read_2_data_T_1377 | _io_read_2_data_T_1363; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_1550 = io_read_2_addr[15] & payload_15_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_1581 = io_read_2_addr[15] & payload_15_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1597 = io_read_2_addr[0] ? payload_0_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1598 = io_read_2_addr[1] ? payload_1_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1599 = io_read_2_addr[2] ? payload_2_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1600 = io_read_2_addr[3] ? payload_3_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1601 = io_read_2_addr[4] ? payload_4_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1602 = io_read_2_addr[5] ? payload_5_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1603 = io_read_2_addr[6] ? payload_6_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1604 = io_read_2_addr[7] ? payload_7_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1605 = io_read_2_addr[8] ? payload_8_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1606 = io_read_2_addr[9] ? payload_9_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1607 = io_read_2_addr[10] ? payload_10_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1608 = io_read_2_addr[11] ? payload_11_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1609 = io_read_2_addr[12] ? payload_12_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1610 = io_read_2_addr[13] ? payload_13_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1611 = io_read_2_addr[14] ? payload_14_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1612 = io_read_2_addr[15] ? payload_15_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1613 = _io_read_2_data_T_1597 | _io_read_2_data_T_1598; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1614 = _io_read_2_data_T_1613 | _io_read_2_data_T_1599; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1615 = _io_read_2_data_T_1614 | _io_read_2_data_T_1600; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1616 = _io_read_2_data_T_1615 | _io_read_2_data_T_1601; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1617 = _io_read_2_data_T_1616 | _io_read_2_data_T_1602; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1618 = _io_read_2_data_T_1617 | _io_read_2_data_T_1603; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1619 = _io_read_2_data_T_1618 | _io_read_2_data_T_1604; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1620 = _io_read_2_data_T_1619 | _io_read_2_data_T_1605; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1621 = _io_read_2_data_T_1620 | _io_read_2_data_T_1606; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1622 = _io_read_2_data_T_1621 | _io_read_2_data_T_1607; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1623 = _io_read_2_data_T_1622 | _io_read_2_data_T_1608; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1624 = _io_read_2_data_T_1623 | _io_read_2_data_T_1609; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1625 = _io_read_2_data_T_1624 | _io_read_2_data_T_1610; // @[Mux.scala 27:73]
  wire [6:0] _io_read_2_data_T_1626 = _io_read_2_data_T_1625 | _io_read_2_data_T_1611; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1628 = io_read_2_addr[0] ? payload_0_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1629 = io_read_2_addr[1] ? payload_1_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1630 = io_read_2_addr[2] ? payload_2_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1631 = io_read_2_addr[3] ? payload_3_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1632 = io_read_2_addr[4] ? payload_4_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1633 = io_read_2_addr[5] ? payload_5_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1634 = io_read_2_addr[6] ? payload_6_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1635 = io_read_2_addr[7] ? payload_7_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1636 = io_read_2_addr[8] ? payload_8_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1637 = io_read_2_addr[9] ? payload_9_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1638 = io_read_2_addr[10] ? payload_10_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1639 = io_read_2_addr[11] ? payload_11_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1640 = io_read_2_addr[12] ? payload_12_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1641 = io_read_2_addr[13] ? payload_13_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1642 = io_read_2_addr[14] ? payload_14_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1643 = io_read_2_addr[15] ? payload_15_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1644 = _io_read_2_data_T_1628 | _io_read_2_data_T_1629; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1645 = _io_read_2_data_T_1644 | _io_read_2_data_T_1630; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1646 = _io_read_2_data_T_1645 | _io_read_2_data_T_1631; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1647 = _io_read_2_data_T_1646 | _io_read_2_data_T_1632; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1648 = _io_read_2_data_T_1647 | _io_read_2_data_T_1633; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1649 = _io_read_2_data_T_1648 | _io_read_2_data_T_1634; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1650 = _io_read_2_data_T_1649 | _io_read_2_data_T_1635; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1651 = _io_read_2_data_T_1650 | _io_read_2_data_T_1636; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1652 = _io_read_2_data_T_1651 | _io_read_2_data_T_1637; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1653 = _io_read_2_data_T_1652 | _io_read_2_data_T_1638; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1654 = _io_read_2_data_T_1653 | _io_read_2_data_T_1639; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1655 = _io_read_2_data_T_1654 | _io_read_2_data_T_1640; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1656 = _io_read_2_data_T_1655 | _io_read_2_data_T_1641; // @[Mux.scala 27:73]
  wire [3:0] _io_read_2_data_T_1657 = _io_read_2_data_T_1656 | _io_read_2_data_T_1642; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1907 = io_read_2_addr[0] ? payload_0_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1908 = io_read_2_addr[1] ? payload_1_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1909 = io_read_2_addr[2] ? payload_2_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1910 = io_read_2_addr[3] ? payload_3_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1911 = io_read_2_addr[4] ? payload_4_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1912 = io_read_2_addr[5] ? payload_5_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1913 = io_read_2_addr[6] ? payload_6_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1914 = io_read_2_addr[7] ? payload_7_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1915 = io_read_2_addr[8] ? payload_8_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1916 = io_read_2_addr[9] ? payload_9_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1917 = io_read_2_addr[10] ? payload_10_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1918 = io_read_2_addr[11] ? payload_11_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1919 = io_read_2_addr[12] ? payload_12_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1920 = io_read_2_addr[13] ? payload_13_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1921 = io_read_2_addr[14] ? payload_14_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1922 = io_read_2_addr[15] ? payload_15_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1923 = _io_read_2_data_T_1907 | _io_read_2_data_T_1908; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1924 = _io_read_2_data_T_1923 | _io_read_2_data_T_1909; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1925 = _io_read_2_data_T_1924 | _io_read_2_data_T_1910; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1926 = _io_read_2_data_T_1925 | _io_read_2_data_T_1911; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1927 = _io_read_2_data_T_1926 | _io_read_2_data_T_1912; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1928 = _io_read_2_data_T_1927 | _io_read_2_data_T_1913; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1929 = _io_read_2_data_T_1928 | _io_read_2_data_T_1914; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1930 = _io_read_2_data_T_1929 | _io_read_2_data_T_1915; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1931 = _io_read_2_data_T_1930 | _io_read_2_data_T_1916; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1932 = _io_read_2_data_T_1931 | _io_read_2_data_T_1917; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1933 = _io_read_2_data_T_1932 | _io_read_2_data_T_1918; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1934 = _io_read_2_data_T_1933 | _io_read_2_data_T_1919; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1935 = _io_read_2_data_T_1934 | _io_read_2_data_T_1920; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1936 = _io_read_2_data_T_1935 | _io_read_2_data_T_1921; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1938 = io_read_2_addr[0] ? payload_0_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1939 = io_read_2_addr[1] ? payload_1_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1940 = io_read_2_addr[2] ? payload_2_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1941 = io_read_2_addr[3] ? payload_3_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1942 = io_read_2_addr[4] ? payload_4_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1943 = io_read_2_addr[5] ? payload_5_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1944 = io_read_2_addr[6] ? payload_6_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1945 = io_read_2_addr[7] ? payload_7_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1946 = io_read_2_addr[8] ? payload_8_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1947 = io_read_2_addr[9] ? payload_9_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1948 = io_read_2_addr[10] ? payload_10_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1949 = io_read_2_addr[11] ? payload_11_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1950 = io_read_2_addr[12] ? payload_12_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1951 = io_read_2_addr[13] ? payload_13_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1952 = io_read_2_addr[14] ? payload_14_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1953 = io_read_2_addr[15] ? payload_15_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1954 = _io_read_2_data_T_1938 | _io_read_2_data_T_1939; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1955 = _io_read_2_data_T_1954 | _io_read_2_data_T_1940; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1956 = _io_read_2_data_T_1955 | _io_read_2_data_T_1941; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1957 = _io_read_2_data_T_1956 | _io_read_2_data_T_1942; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1958 = _io_read_2_data_T_1957 | _io_read_2_data_T_1943; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1959 = _io_read_2_data_T_1958 | _io_read_2_data_T_1944; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1960 = _io_read_2_data_T_1959 | _io_read_2_data_T_1945; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1961 = _io_read_2_data_T_1960 | _io_read_2_data_T_1946; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1962 = _io_read_2_data_T_1961 | _io_read_2_data_T_1947; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1963 = _io_read_2_data_T_1962 | _io_read_2_data_T_1948; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1964 = _io_read_2_data_T_1963 | _io_read_2_data_T_1949; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1965 = _io_read_2_data_T_1964 | _io_read_2_data_T_1950; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1966 = _io_read_2_data_T_1965 | _io_read_2_data_T_1951; // @[Mux.scala 27:73]
  wire [2:0] _io_read_2_data_T_1967 = _io_read_2_data_T_1966 | _io_read_2_data_T_1952; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_1984 = io_read_2_addr[15] & payload_15_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2000 = io_read_2_addr[0] ? payload_0_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2001 = io_read_2_addr[1] ? payload_1_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2002 = io_read_2_addr[2] ? payload_2_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2003 = io_read_2_addr[3] ? payload_3_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2004 = io_read_2_addr[4] ? payload_4_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2005 = io_read_2_addr[5] ? payload_5_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2006 = io_read_2_addr[6] ? payload_6_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2007 = io_read_2_addr[7] ? payload_7_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2008 = io_read_2_addr[8] ? payload_8_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2009 = io_read_2_addr[9] ? payload_9_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2010 = io_read_2_addr[10] ? payload_10_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2011 = io_read_2_addr[11] ? payload_11_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2012 = io_read_2_addr[12] ? payload_12_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2013 = io_read_2_addr[13] ? payload_13_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2014 = io_read_2_addr[14] ? payload_14_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2015 = io_read_2_addr[15] ? payload_15_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2016 = _io_read_2_data_T_2000 | _io_read_2_data_T_2001; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2017 = _io_read_2_data_T_2016 | _io_read_2_data_T_2002; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2018 = _io_read_2_data_T_2017 | _io_read_2_data_T_2003; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2019 = _io_read_2_data_T_2018 | _io_read_2_data_T_2004; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2020 = _io_read_2_data_T_2019 | _io_read_2_data_T_2005; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2021 = _io_read_2_data_T_2020 | _io_read_2_data_T_2006; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2022 = _io_read_2_data_T_2021 | _io_read_2_data_T_2007; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2023 = _io_read_2_data_T_2022 | _io_read_2_data_T_2008; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2024 = _io_read_2_data_T_2023 | _io_read_2_data_T_2009; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2025 = _io_read_2_data_T_2024 | _io_read_2_data_T_2010; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2026 = _io_read_2_data_T_2025 | _io_read_2_data_T_2011; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2027 = _io_read_2_data_T_2026 | _io_read_2_data_T_2012; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2028 = _io_read_2_data_T_2027 | _io_read_2_data_T_2013; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2029 = _io_read_2_data_T_2028 | _io_read_2_data_T_2014; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2046 = io_read_2_addr[15] & payload_15_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2077 = io_read_2_addr[15] & payload_15_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2093 = io_read_2_addr[0] ? payload_0_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2094 = io_read_2_addr[1] ? payload_1_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2095 = io_read_2_addr[2] ? payload_2_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2096 = io_read_2_addr[3] ? payload_3_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2097 = io_read_2_addr[4] ? payload_4_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2098 = io_read_2_addr[5] ? payload_5_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2099 = io_read_2_addr[6] ? payload_6_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2100 = io_read_2_addr[7] ? payload_7_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2101 = io_read_2_addr[8] ? payload_8_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2102 = io_read_2_addr[9] ? payload_9_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2103 = io_read_2_addr[10] ? payload_10_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2104 = io_read_2_addr[11] ? payload_11_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2105 = io_read_2_addr[12] ? payload_12_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2106 = io_read_2_addr[13] ? payload_13_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2107 = io_read_2_addr[14] ? payload_14_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2108 = io_read_2_addr[15] ? payload_15_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2109 = _io_read_2_data_T_2093 | _io_read_2_data_T_2094; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2110 = _io_read_2_data_T_2109 | _io_read_2_data_T_2095; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2111 = _io_read_2_data_T_2110 | _io_read_2_data_T_2096; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2112 = _io_read_2_data_T_2111 | _io_read_2_data_T_2097; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2113 = _io_read_2_data_T_2112 | _io_read_2_data_T_2098; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2114 = _io_read_2_data_T_2113 | _io_read_2_data_T_2099; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2115 = _io_read_2_data_T_2114 | _io_read_2_data_T_2100; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2116 = _io_read_2_data_T_2115 | _io_read_2_data_T_2101; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2117 = _io_read_2_data_T_2116 | _io_read_2_data_T_2102; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2118 = _io_read_2_data_T_2117 | _io_read_2_data_T_2103; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2119 = _io_read_2_data_T_2118 | _io_read_2_data_T_2104; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2120 = _io_read_2_data_T_2119 | _io_read_2_data_T_2105; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2121 = _io_read_2_data_T_2120 | _io_read_2_data_T_2106; // @[Mux.scala 27:73]
  wire [4:0] _io_read_2_data_T_2122 = _io_read_2_data_T_2121 | _io_read_2_data_T_2107; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2139 = io_read_2_addr[15] & payload_15_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2170 = io_read_2_addr[15] & payload_15_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2232 = io_read_2_addr[15] & payload_15_cf_pred_taken; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2263 = io_read_2_addr[15] & payload_15_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2294 = io_read_2_addr[15] & payload_15_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2310 = io_read_2_addr[0] ? payload_0_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2311 = io_read_2_addr[1] ? payload_1_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2312 = io_read_2_addr[2] ? payload_2_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2313 = io_read_2_addr[3] ? payload_3_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2314 = io_read_2_addr[4] ? payload_4_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2315 = io_read_2_addr[5] ? payload_5_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2316 = io_read_2_addr[6] ? payload_6_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2317 = io_read_2_addr[7] ? payload_7_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2318 = io_read_2_addr[8] ? payload_8_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2319 = io_read_2_addr[9] ? payload_9_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2320 = io_read_2_addr[10] ? payload_10_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2321 = io_read_2_addr[11] ? payload_11_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2322 = io_read_2_addr[12] ? payload_12_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2323 = io_read_2_addr[13] ? payload_13_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2324 = io_read_2_addr[14] ? payload_14_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2325 = io_read_2_addr[15] ? payload_15_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2326 = _io_read_2_data_T_2310 | _io_read_2_data_T_2311; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2327 = _io_read_2_data_T_2326 | _io_read_2_data_T_2312; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2328 = _io_read_2_data_T_2327 | _io_read_2_data_T_2313; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2329 = _io_read_2_data_T_2328 | _io_read_2_data_T_2314; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2330 = _io_read_2_data_T_2329 | _io_read_2_data_T_2315; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2331 = _io_read_2_data_T_2330 | _io_read_2_data_T_2316; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2332 = _io_read_2_data_T_2331 | _io_read_2_data_T_2317; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2333 = _io_read_2_data_T_2332 | _io_read_2_data_T_2318; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2334 = _io_read_2_data_T_2333 | _io_read_2_data_T_2319; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2335 = _io_read_2_data_T_2334 | _io_read_2_data_T_2320; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2336 = _io_read_2_data_T_2335 | _io_read_2_data_T_2321; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2337 = _io_read_2_data_T_2336 | _io_read_2_data_T_2322; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2338 = _io_read_2_data_T_2337 | _io_read_2_data_T_2323; // @[Mux.scala 27:73]
  wire [1:0] _io_read_2_data_T_2339 = _io_read_2_data_T_2338 | _io_read_2_data_T_2324; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2356 = io_read_2_addr[15] & payload_15_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2604 = io_read_2_addr[15] & payload_15_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  _io_read_2_data_T_2635 = io_read_2_addr[15] & payload_15_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3271 = io_read_2_addr[0] ? payload_0_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3272 = io_read_2_addr[1] ? payload_1_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3273 = io_read_2_addr[2] ? payload_2_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3274 = io_read_2_addr[3] ? payload_3_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3275 = io_read_2_addr[4] ? payload_4_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3276 = io_read_2_addr[5] ? payload_5_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3277 = io_read_2_addr[6] ? payload_6_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3278 = io_read_2_addr[7] ? payload_7_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3279 = io_read_2_addr[8] ? payload_8_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3280 = io_read_2_addr[9] ? payload_9_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3281 = io_read_2_addr[10] ? payload_10_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3282 = io_read_2_addr[11] ? payload_11_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3283 = io_read_2_addr[12] ? payload_12_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3284 = io_read_2_addr[13] ? payload_13_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3285 = io_read_2_addr[14] ? payload_14_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3286 = io_read_2_addr[15] ? payload_15_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3287 = _io_read_2_data_T_3271 | _io_read_2_data_T_3272; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3288 = _io_read_2_data_T_3287 | _io_read_2_data_T_3273; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3289 = _io_read_2_data_T_3288 | _io_read_2_data_T_3274; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3290 = _io_read_2_data_T_3289 | _io_read_2_data_T_3275; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3291 = _io_read_2_data_T_3290 | _io_read_2_data_T_3276; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3292 = _io_read_2_data_T_3291 | _io_read_2_data_T_3277; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3293 = _io_read_2_data_T_3292 | _io_read_2_data_T_3278; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3294 = _io_read_2_data_T_3293 | _io_read_2_data_T_3279; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3295 = _io_read_2_data_T_3294 | _io_read_2_data_T_3280; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3296 = _io_read_2_data_T_3295 | _io_read_2_data_T_3281; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3297 = _io_read_2_data_T_3296 | _io_read_2_data_T_3282; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3298 = _io_read_2_data_T_3297 | _io_read_2_data_T_3283; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3299 = _io_read_2_data_T_3298 | _io_read_2_data_T_3284; // @[Mux.scala 27:73]
  wire [9:0] _io_read_2_data_T_3300 = _io_read_2_data_T_3299 | _io_read_2_data_T_3285; // @[Mux.scala 27:73]
  wire  wenVec__0 = io_write_0_enable & io_write_0_addr[0]; // @[PayloadArray.scala 55:53]
  wire  wenVec__1 = io_write_1_enable & io_write_1_addr[0]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T = {wenVec__1,wenVec__0}; // @[PayloadArray.scala 56:22]
  wire  wen = |_wen_T; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_33 = wenVec__0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_34 = wenVec__1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_sqIdx_value = _wdata_T_33 | _wdata_T_34; // @[Mux.scala 27:73]
  wire  wdata_sqIdx_flag = wenVec__0 & io_write_0_data_sqIdx_flag | wenVec__1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_39 = wenVec__0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_40 = wenVec__1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_lqIdx_value = _wdata_T_39 | _wdata_T_40; // @[Mux.scala 27:73]
  wire  wdata_lqIdx_flag = wenVec__0 & io_write_0_data_lqIdx_flag | wenVec__1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_45 = wenVec__0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_46 = wenVec__1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_robIdx_value = _wdata_T_45 | _wdata_T_46; // @[Mux.scala 27:73]
  wire  wdata_robIdx_flag = wenVec__0 & io_write_0_data_robIdx_flag | wenVec__1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_54 = wenVec__0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_55 = wenVec__1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_pdest = _wdata_T_54 | _wdata_T_55; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_129 = wenVec__0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_130 = wenVec__1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_ctrl_imm = _wdata_T_129 | _wdata_T_130; // @[Mux.scala 27:73]
  wire  wdata_ctrl_fpWen = wenVec__0 & io_write_0_data_ctrl_fpWen | wenVec__1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_ctrl_rfWen = wenVec__0 & io_write_0_data_ctrl_rfWen | wenVec__1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_153 = wenVec__0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_154 = wenVec__1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_ctrl_fuOpType = _wdata_T_153 | _wdata_T_154; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_156 = wenVec__0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_157 = wenVec__1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_ctrl_fuType = _wdata_T_156 | _wdata_T_157; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_183 = wenVec__0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_184 = wenVec__1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_cf_ftqOffset = _wdata_T_183 | _wdata_T_184; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_186 = wenVec__0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_187 = wenVec__1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_cf_ftqPtr_value = _wdata_T_186 | _wdata_T_187; // @[Mux.scala 27:73]
  wire  wdata_cf_ftqPtr_flag = wenVec__0 & io_write_0_data_cf_ftqPtr_flag | wenVec__1 & io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_192 = wenVec__0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_193 = wenVec__1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_cf_ssid = _wdata_T_192 | _wdata_T_193; // @[Mux.scala 27:73]
  wire  wdata_cf_loadWaitStrict = wenVec__0 & io_write_0_data_cf_loadWaitStrict | wenVec__1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_cf_loadWaitBit = wenVec__0 & io_write_0_data_cf_loadWaitBit | wenVec__1 & io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_201 = wenVec__0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_202 = wenVec__1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_cf_waitForRobIdx_value = _wdata_T_201 | _wdata_T_202; // @[Mux.scala 27:73]
  wire  wdata_cf_waitForRobIdx_flag = wenVec__0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec__1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_cf_storeSetHit = wenVec__0 & io_write_0_data_cf_storeSetHit | wenVec__1 & io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_cf_pred_taken = wenVec__0 & io_write_0_data_cf_pred_taken | wenVec__1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_cf_pd_isRet = wenVec__0 & io_write_0_data_cf_pd_isRet | wenVec__1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_cf_pd_isCall = wenVec__0 & io_write_0_data_cf_pd_isCall | wenVec__1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_222 = wenVec__0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_223 = wenVec__1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_cf_pd_brType = _wdata_T_222 | _wdata_T_223; // @[Mux.scala 27:73]
  wire  wdata_cf_pd_isRVC = wenVec__0 & io_write_0_data_cf_pd_isRVC | wenVec__1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_cf_trigger_backendEn_0 = wenVec__0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec__1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_cf_trigger_backendEn_1 = wenVec__0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec__1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_315 = wenVec__0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_316 = wenVec__1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_cf_foldpc = _wdata_T_315 | _wdata_T_316; // @[Mux.scala 27:73]
  wire  wenVec_1_0 = io_write_0_enable & io_write_0_addr[1]; // @[PayloadArray.scala 55:53]
  wire  wenVec_1_1 = io_write_1_enable & io_write_1_addr[1]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_1 = {wenVec_1_1,wenVec_1_0}; // @[PayloadArray.scala 56:22]
  wire  wen_1 = |_wen_T_1; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_357 = wenVec_1_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_358 = wenVec_1_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_1_sqIdx_value = _wdata_T_357 | _wdata_T_358; // @[Mux.scala 27:73]
  wire  wdata_1_sqIdx_flag = wenVec_1_0 & io_write_0_data_sqIdx_flag | wenVec_1_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_363 = wenVec_1_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_364 = wenVec_1_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_1_lqIdx_value = _wdata_T_363 | _wdata_T_364; // @[Mux.scala 27:73]
  wire  wdata_1_lqIdx_flag = wenVec_1_0 & io_write_0_data_lqIdx_flag | wenVec_1_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_369 = wenVec_1_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_370 = wenVec_1_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_1_robIdx_value = _wdata_T_369 | _wdata_T_370; // @[Mux.scala 27:73]
  wire  wdata_1_robIdx_flag = wenVec_1_0 & io_write_0_data_robIdx_flag | wenVec_1_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_378 = wenVec_1_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_379 = wenVec_1_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_1_pdest = _wdata_T_378 | _wdata_T_379; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_453 = wenVec_1_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_454 = wenVec_1_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_1_ctrl_imm = _wdata_T_453 | _wdata_T_454; // @[Mux.scala 27:73]
  wire  wdata_1_ctrl_fpWen = wenVec_1_0 & io_write_0_data_ctrl_fpWen | wenVec_1_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_1_ctrl_rfWen = wenVec_1_0 & io_write_0_data_ctrl_rfWen | wenVec_1_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_477 = wenVec_1_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_478 = wenVec_1_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_1_ctrl_fuOpType = _wdata_T_477 | _wdata_T_478; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_480 = wenVec_1_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_481 = wenVec_1_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_1_ctrl_fuType = _wdata_T_480 | _wdata_T_481; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_507 = wenVec_1_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_508 = wenVec_1_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_1_cf_ftqOffset = _wdata_T_507 | _wdata_T_508; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_510 = wenVec_1_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_511 = wenVec_1_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_1_cf_ftqPtr_value = _wdata_T_510 | _wdata_T_511; // @[Mux.scala 27:73]
  wire  wdata_1_cf_ftqPtr_flag = wenVec_1_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_1_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_516 = wenVec_1_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_517 = wenVec_1_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_1_cf_ssid = _wdata_T_516 | _wdata_T_517; // @[Mux.scala 27:73]
  wire  wdata_1_cf_loadWaitStrict = wenVec_1_0 & io_write_0_data_cf_loadWaitStrict | wenVec_1_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_1_cf_loadWaitBit = wenVec_1_0 & io_write_0_data_cf_loadWaitBit | wenVec_1_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_525 = wenVec_1_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_526 = wenVec_1_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_1_cf_waitForRobIdx_value = _wdata_T_525 | _wdata_T_526; // @[Mux.scala 27:73]
  wire  wdata_1_cf_waitForRobIdx_flag = wenVec_1_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_1_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_1_cf_storeSetHit = wenVec_1_0 & io_write_0_data_cf_storeSetHit | wenVec_1_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_1_cf_pred_taken = wenVec_1_0 & io_write_0_data_cf_pred_taken | wenVec_1_1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_1_cf_pd_isRet = wenVec_1_0 & io_write_0_data_cf_pd_isRet | wenVec_1_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_1_cf_pd_isCall = wenVec_1_0 & io_write_0_data_cf_pd_isCall | wenVec_1_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_546 = wenVec_1_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_547 = wenVec_1_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_1_cf_pd_brType = _wdata_T_546 | _wdata_T_547; // @[Mux.scala 27:73]
  wire  wdata_1_cf_pd_isRVC = wenVec_1_0 & io_write_0_data_cf_pd_isRVC | wenVec_1_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_1_cf_trigger_backendEn_0 = wenVec_1_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_1_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_1_cf_trigger_backendEn_1 = wenVec_1_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_1_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_639 = wenVec_1_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_640 = wenVec_1_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_1_cf_foldpc = _wdata_T_639 | _wdata_T_640; // @[Mux.scala 27:73]
  wire  wenVec_2_0 = io_write_0_enable & io_write_0_addr[2]; // @[PayloadArray.scala 55:53]
  wire  wenVec_2_1 = io_write_1_enable & io_write_1_addr[2]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_2 = {wenVec_2_1,wenVec_2_0}; // @[PayloadArray.scala 56:22]
  wire  wen_2 = |_wen_T_2; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_681 = wenVec_2_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_682 = wenVec_2_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_2_sqIdx_value = _wdata_T_681 | _wdata_T_682; // @[Mux.scala 27:73]
  wire  wdata_2_sqIdx_flag = wenVec_2_0 & io_write_0_data_sqIdx_flag | wenVec_2_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_687 = wenVec_2_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_688 = wenVec_2_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_2_lqIdx_value = _wdata_T_687 | _wdata_T_688; // @[Mux.scala 27:73]
  wire  wdata_2_lqIdx_flag = wenVec_2_0 & io_write_0_data_lqIdx_flag | wenVec_2_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_693 = wenVec_2_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_694 = wenVec_2_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_2_robIdx_value = _wdata_T_693 | _wdata_T_694; // @[Mux.scala 27:73]
  wire  wdata_2_robIdx_flag = wenVec_2_0 & io_write_0_data_robIdx_flag | wenVec_2_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_702 = wenVec_2_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_703 = wenVec_2_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_2_pdest = _wdata_T_702 | _wdata_T_703; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_777 = wenVec_2_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_778 = wenVec_2_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_2_ctrl_imm = _wdata_T_777 | _wdata_T_778; // @[Mux.scala 27:73]
  wire  wdata_2_ctrl_fpWen = wenVec_2_0 & io_write_0_data_ctrl_fpWen | wenVec_2_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_2_ctrl_rfWen = wenVec_2_0 & io_write_0_data_ctrl_rfWen | wenVec_2_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_801 = wenVec_2_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_802 = wenVec_2_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_2_ctrl_fuOpType = _wdata_T_801 | _wdata_T_802; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_804 = wenVec_2_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_805 = wenVec_2_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_2_ctrl_fuType = _wdata_T_804 | _wdata_T_805; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_831 = wenVec_2_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_832 = wenVec_2_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_2_cf_ftqOffset = _wdata_T_831 | _wdata_T_832; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_834 = wenVec_2_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_835 = wenVec_2_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_2_cf_ftqPtr_value = _wdata_T_834 | _wdata_T_835; // @[Mux.scala 27:73]
  wire  wdata_2_cf_ftqPtr_flag = wenVec_2_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_2_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_840 = wenVec_2_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_841 = wenVec_2_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_2_cf_ssid = _wdata_T_840 | _wdata_T_841; // @[Mux.scala 27:73]
  wire  wdata_2_cf_loadWaitStrict = wenVec_2_0 & io_write_0_data_cf_loadWaitStrict | wenVec_2_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_2_cf_loadWaitBit = wenVec_2_0 & io_write_0_data_cf_loadWaitBit | wenVec_2_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_849 = wenVec_2_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_850 = wenVec_2_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_2_cf_waitForRobIdx_value = _wdata_T_849 | _wdata_T_850; // @[Mux.scala 27:73]
  wire  wdata_2_cf_waitForRobIdx_flag = wenVec_2_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_2_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_2_cf_storeSetHit = wenVec_2_0 & io_write_0_data_cf_storeSetHit | wenVec_2_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_2_cf_pred_taken = wenVec_2_0 & io_write_0_data_cf_pred_taken | wenVec_2_1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_2_cf_pd_isRet = wenVec_2_0 & io_write_0_data_cf_pd_isRet | wenVec_2_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_2_cf_pd_isCall = wenVec_2_0 & io_write_0_data_cf_pd_isCall | wenVec_2_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_870 = wenVec_2_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_871 = wenVec_2_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_2_cf_pd_brType = _wdata_T_870 | _wdata_T_871; // @[Mux.scala 27:73]
  wire  wdata_2_cf_pd_isRVC = wenVec_2_0 & io_write_0_data_cf_pd_isRVC | wenVec_2_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_2_cf_trigger_backendEn_0 = wenVec_2_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_2_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_2_cf_trigger_backendEn_1 = wenVec_2_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_2_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_963 = wenVec_2_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_964 = wenVec_2_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_2_cf_foldpc = _wdata_T_963 | _wdata_T_964; // @[Mux.scala 27:73]
  wire  wenVec_3_0 = io_write_0_enable & io_write_0_addr[3]; // @[PayloadArray.scala 55:53]
  wire  wenVec_3_1 = io_write_1_enable & io_write_1_addr[3]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_3 = {wenVec_3_1,wenVec_3_0}; // @[PayloadArray.scala 56:22]
  wire  wen_3 = |_wen_T_3; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_1005 = wenVec_3_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1006 = wenVec_3_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_3_sqIdx_value = _wdata_T_1005 | _wdata_T_1006; // @[Mux.scala 27:73]
  wire  wdata_3_sqIdx_flag = wenVec_3_0 & io_write_0_data_sqIdx_flag | wenVec_3_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1011 = wenVec_3_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1012 = wenVec_3_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_3_lqIdx_value = _wdata_T_1011 | _wdata_T_1012; // @[Mux.scala 27:73]
  wire  wdata_3_lqIdx_flag = wenVec_3_0 & io_write_0_data_lqIdx_flag | wenVec_3_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1017 = wenVec_3_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1018 = wenVec_3_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_3_robIdx_value = _wdata_T_1017 | _wdata_T_1018; // @[Mux.scala 27:73]
  wire  wdata_3_robIdx_flag = wenVec_3_0 & io_write_0_data_robIdx_flag | wenVec_3_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_1026 = wenVec_3_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_1027 = wenVec_3_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_3_pdest = _wdata_T_1026 | _wdata_T_1027; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_1101 = wenVec_3_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_1102 = wenVec_3_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_3_ctrl_imm = _wdata_T_1101 | _wdata_T_1102; // @[Mux.scala 27:73]
  wire  wdata_3_ctrl_fpWen = wenVec_3_0 & io_write_0_data_ctrl_fpWen | wenVec_3_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_3_ctrl_rfWen = wenVec_3_0 & io_write_0_data_ctrl_rfWen | wenVec_3_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_1125 = wenVec_3_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_1126 = wenVec_3_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_3_ctrl_fuOpType = _wdata_T_1125 | _wdata_T_1126; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1128 = wenVec_3_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1129 = wenVec_3_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_3_ctrl_fuType = _wdata_T_1128 | _wdata_T_1129; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1155 = wenVec_3_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1156 = wenVec_3_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_3_cf_ftqOffset = _wdata_T_1155 | _wdata_T_1156; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1158 = wenVec_3_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1159 = wenVec_3_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_3_cf_ftqPtr_value = _wdata_T_1158 | _wdata_T_1159; // @[Mux.scala 27:73]
  wire  wdata_3_cf_ftqPtr_flag = wenVec_3_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_3_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1164 = wenVec_3_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1165 = wenVec_3_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_3_cf_ssid = _wdata_T_1164 | _wdata_T_1165; // @[Mux.scala 27:73]
  wire  wdata_3_cf_loadWaitStrict = wenVec_3_0 & io_write_0_data_cf_loadWaitStrict | wenVec_3_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_3_cf_loadWaitBit = wenVec_3_0 & io_write_0_data_cf_loadWaitBit | wenVec_3_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1173 = wenVec_3_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1174 = wenVec_3_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_3_cf_waitForRobIdx_value = _wdata_T_1173 | _wdata_T_1174; // @[Mux.scala 27:73]
  wire  wdata_3_cf_waitForRobIdx_flag = wenVec_3_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_3_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_3_cf_storeSetHit = wenVec_3_0 & io_write_0_data_cf_storeSetHit | wenVec_3_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_3_cf_pred_taken = wenVec_3_0 & io_write_0_data_cf_pred_taken | wenVec_3_1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_3_cf_pd_isRet = wenVec_3_0 & io_write_0_data_cf_pd_isRet | wenVec_3_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_3_cf_pd_isCall = wenVec_3_0 & io_write_0_data_cf_pd_isCall | wenVec_3_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_1194 = wenVec_3_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_1195 = wenVec_3_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_3_cf_pd_brType = _wdata_T_1194 | _wdata_T_1195; // @[Mux.scala 27:73]
  wire  wdata_3_cf_pd_isRVC = wenVec_3_0 & io_write_0_data_cf_pd_isRVC | wenVec_3_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_3_cf_trigger_backendEn_0 = wenVec_3_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_3_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_3_cf_trigger_backendEn_1 = wenVec_3_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_3_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_1287 = wenVec_3_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_1288 = wenVec_3_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_3_cf_foldpc = _wdata_T_1287 | _wdata_T_1288; // @[Mux.scala 27:73]
  wire  wenVec_4_0 = io_write_0_enable & io_write_0_addr[4]; // @[PayloadArray.scala 55:53]
  wire  wenVec_4_1 = io_write_1_enable & io_write_1_addr[4]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_4 = {wenVec_4_1,wenVec_4_0}; // @[PayloadArray.scala 56:22]
  wire  wen_4 = |_wen_T_4; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_1329 = wenVec_4_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1330 = wenVec_4_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_4_sqIdx_value = _wdata_T_1329 | _wdata_T_1330; // @[Mux.scala 27:73]
  wire  wdata_4_sqIdx_flag = wenVec_4_0 & io_write_0_data_sqIdx_flag | wenVec_4_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1335 = wenVec_4_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1336 = wenVec_4_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_4_lqIdx_value = _wdata_T_1335 | _wdata_T_1336; // @[Mux.scala 27:73]
  wire  wdata_4_lqIdx_flag = wenVec_4_0 & io_write_0_data_lqIdx_flag | wenVec_4_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1341 = wenVec_4_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1342 = wenVec_4_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_4_robIdx_value = _wdata_T_1341 | _wdata_T_1342; // @[Mux.scala 27:73]
  wire  wdata_4_robIdx_flag = wenVec_4_0 & io_write_0_data_robIdx_flag | wenVec_4_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_1350 = wenVec_4_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_1351 = wenVec_4_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_4_pdest = _wdata_T_1350 | _wdata_T_1351; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_1425 = wenVec_4_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_1426 = wenVec_4_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_4_ctrl_imm = _wdata_T_1425 | _wdata_T_1426; // @[Mux.scala 27:73]
  wire  wdata_4_ctrl_fpWen = wenVec_4_0 & io_write_0_data_ctrl_fpWen | wenVec_4_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_4_ctrl_rfWen = wenVec_4_0 & io_write_0_data_ctrl_rfWen | wenVec_4_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_1449 = wenVec_4_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_1450 = wenVec_4_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_4_ctrl_fuOpType = _wdata_T_1449 | _wdata_T_1450; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1452 = wenVec_4_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1453 = wenVec_4_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_4_ctrl_fuType = _wdata_T_1452 | _wdata_T_1453; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1479 = wenVec_4_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1480 = wenVec_4_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_4_cf_ftqOffset = _wdata_T_1479 | _wdata_T_1480; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1482 = wenVec_4_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1483 = wenVec_4_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_4_cf_ftqPtr_value = _wdata_T_1482 | _wdata_T_1483; // @[Mux.scala 27:73]
  wire  wdata_4_cf_ftqPtr_flag = wenVec_4_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_4_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1488 = wenVec_4_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1489 = wenVec_4_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_4_cf_ssid = _wdata_T_1488 | _wdata_T_1489; // @[Mux.scala 27:73]
  wire  wdata_4_cf_loadWaitStrict = wenVec_4_0 & io_write_0_data_cf_loadWaitStrict | wenVec_4_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_4_cf_loadWaitBit = wenVec_4_0 & io_write_0_data_cf_loadWaitBit | wenVec_4_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1497 = wenVec_4_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1498 = wenVec_4_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_4_cf_waitForRobIdx_value = _wdata_T_1497 | _wdata_T_1498; // @[Mux.scala 27:73]
  wire  wdata_4_cf_waitForRobIdx_flag = wenVec_4_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_4_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_4_cf_storeSetHit = wenVec_4_0 & io_write_0_data_cf_storeSetHit | wenVec_4_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_4_cf_pred_taken = wenVec_4_0 & io_write_0_data_cf_pred_taken | wenVec_4_1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_4_cf_pd_isRet = wenVec_4_0 & io_write_0_data_cf_pd_isRet | wenVec_4_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_4_cf_pd_isCall = wenVec_4_0 & io_write_0_data_cf_pd_isCall | wenVec_4_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_1518 = wenVec_4_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_1519 = wenVec_4_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_4_cf_pd_brType = _wdata_T_1518 | _wdata_T_1519; // @[Mux.scala 27:73]
  wire  wdata_4_cf_pd_isRVC = wenVec_4_0 & io_write_0_data_cf_pd_isRVC | wenVec_4_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_4_cf_trigger_backendEn_0 = wenVec_4_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_4_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_4_cf_trigger_backendEn_1 = wenVec_4_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_4_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_1611 = wenVec_4_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_1612 = wenVec_4_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_4_cf_foldpc = _wdata_T_1611 | _wdata_T_1612; // @[Mux.scala 27:73]
  wire  wenVec_5_0 = io_write_0_enable & io_write_0_addr[5]; // @[PayloadArray.scala 55:53]
  wire  wenVec_5_1 = io_write_1_enable & io_write_1_addr[5]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_5 = {wenVec_5_1,wenVec_5_0}; // @[PayloadArray.scala 56:22]
  wire  wen_5 = |_wen_T_5; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_1653 = wenVec_5_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1654 = wenVec_5_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_5_sqIdx_value = _wdata_T_1653 | _wdata_T_1654; // @[Mux.scala 27:73]
  wire  wdata_5_sqIdx_flag = wenVec_5_0 & io_write_0_data_sqIdx_flag | wenVec_5_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1659 = wenVec_5_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1660 = wenVec_5_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_5_lqIdx_value = _wdata_T_1659 | _wdata_T_1660; // @[Mux.scala 27:73]
  wire  wdata_5_lqIdx_flag = wenVec_5_0 & io_write_0_data_lqIdx_flag | wenVec_5_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1665 = wenVec_5_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1666 = wenVec_5_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_5_robIdx_value = _wdata_T_1665 | _wdata_T_1666; // @[Mux.scala 27:73]
  wire  wdata_5_robIdx_flag = wenVec_5_0 & io_write_0_data_robIdx_flag | wenVec_5_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_1674 = wenVec_5_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_1675 = wenVec_5_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_5_pdest = _wdata_T_1674 | _wdata_T_1675; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_1749 = wenVec_5_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_1750 = wenVec_5_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_5_ctrl_imm = _wdata_T_1749 | _wdata_T_1750; // @[Mux.scala 27:73]
  wire  wdata_5_ctrl_fpWen = wenVec_5_0 & io_write_0_data_ctrl_fpWen | wenVec_5_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_5_ctrl_rfWen = wenVec_5_0 & io_write_0_data_ctrl_rfWen | wenVec_5_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_1773 = wenVec_5_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_1774 = wenVec_5_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_5_ctrl_fuOpType = _wdata_T_1773 | _wdata_T_1774; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1776 = wenVec_5_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1777 = wenVec_5_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_5_ctrl_fuType = _wdata_T_1776 | _wdata_T_1777; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1803 = wenVec_5_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1804 = wenVec_5_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_5_cf_ftqOffset = _wdata_T_1803 | _wdata_T_1804; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1806 = wenVec_5_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_1807 = wenVec_5_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_5_cf_ftqPtr_value = _wdata_T_1806 | _wdata_T_1807; // @[Mux.scala 27:73]
  wire  wdata_5_cf_ftqPtr_flag = wenVec_5_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_5_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1812 = wenVec_5_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1813 = wenVec_5_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_5_cf_ssid = _wdata_T_1812 | _wdata_T_1813; // @[Mux.scala 27:73]
  wire  wdata_5_cf_loadWaitStrict = wenVec_5_0 & io_write_0_data_cf_loadWaitStrict | wenVec_5_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_5_cf_loadWaitBit = wenVec_5_0 & io_write_0_data_cf_loadWaitBit | wenVec_5_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1821 = wenVec_5_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1822 = wenVec_5_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_5_cf_waitForRobIdx_value = _wdata_T_1821 | _wdata_T_1822; // @[Mux.scala 27:73]
  wire  wdata_5_cf_waitForRobIdx_flag = wenVec_5_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_5_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_5_cf_storeSetHit = wenVec_5_0 & io_write_0_data_cf_storeSetHit | wenVec_5_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_5_cf_pred_taken = wenVec_5_0 & io_write_0_data_cf_pred_taken | wenVec_5_1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_5_cf_pd_isRet = wenVec_5_0 & io_write_0_data_cf_pd_isRet | wenVec_5_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_5_cf_pd_isCall = wenVec_5_0 & io_write_0_data_cf_pd_isCall | wenVec_5_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_1842 = wenVec_5_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_1843 = wenVec_5_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_5_cf_pd_brType = _wdata_T_1842 | _wdata_T_1843; // @[Mux.scala 27:73]
  wire  wdata_5_cf_pd_isRVC = wenVec_5_0 & io_write_0_data_cf_pd_isRVC | wenVec_5_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_5_cf_trigger_backendEn_0 = wenVec_5_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_5_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_5_cf_trigger_backendEn_1 = wenVec_5_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_5_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_1935 = wenVec_5_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_1936 = wenVec_5_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_5_cf_foldpc = _wdata_T_1935 | _wdata_T_1936; // @[Mux.scala 27:73]
  wire  wenVec_6_0 = io_write_0_enable & io_write_0_addr[6]; // @[PayloadArray.scala 55:53]
  wire  wenVec_6_1 = io_write_1_enable & io_write_1_addr[6]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_6 = {wenVec_6_1,wenVec_6_0}; // @[PayloadArray.scala 56:22]
  wire  wen_6 = |_wen_T_6; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_1977 = wenVec_6_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1978 = wenVec_6_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_6_sqIdx_value = _wdata_T_1977 | _wdata_T_1978; // @[Mux.scala 27:73]
  wire  wdata_6_sqIdx_flag = wenVec_6_0 & io_write_0_data_sqIdx_flag | wenVec_6_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1983 = wenVec_6_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_1984 = wenVec_6_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_6_lqIdx_value = _wdata_T_1983 | _wdata_T_1984; // @[Mux.scala 27:73]
  wire  wdata_6_lqIdx_flag = wenVec_6_0 & io_write_0_data_lqIdx_flag | wenVec_6_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1989 = wenVec_6_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_1990 = wenVec_6_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_6_robIdx_value = _wdata_T_1989 | _wdata_T_1990; // @[Mux.scala 27:73]
  wire  wdata_6_robIdx_flag = wenVec_6_0 & io_write_0_data_robIdx_flag | wenVec_6_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_1998 = wenVec_6_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_1999 = wenVec_6_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_6_pdest = _wdata_T_1998 | _wdata_T_1999; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_2073 = wenVec_6_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_2074 = wenVec_6_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_6_ctrl_imm = _wdata_T_2073 | _wdata_T_2074; // @[Mux.scala 27:73]
  wire  wdata_6_ctrl_fpWen = wenVec_6_0 & io_write_0_data_ctrl_fpWen | wenVec_6_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_6_ctrl_rfWen = wenVec_6_0 & io_write_0_data_ctrl_rfWen | wenVec_6_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_2097 = wenVec_6_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_2098 = wenVec_6_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_6_ctrl_fuOpType = _wdata_T_2097 | _wdata_T_2098; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2100 = wenVec_6_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2101 = wenVec_6_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_6_ctrl_fuType = _wdata_T_2100 | _wdata_T_2101; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2127 = wenVec_6_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2128 = wenVec_6_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_6_cf_ftqOffset = _wdata_T_2127 | _wdata_T_2128; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2130 = wenVec_6_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2131 = wenVec_6_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_6_cf_ftqPtr_value = _wdata_T_2130 | _wdata_T_2131; // @[Mux.scala 27:73]
  wire  wdata_6_cf_ftqPtr_flag = wenVec_6_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_6_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2136 = wenVec_6_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2137 = wenVec_6_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_6_cf_ssid = _wdata_T_2136 | _wdata_T_2137; // @[Mux.scala 27:73]
  wire  wdata_6_cf_loadWaitStrict = wenVec_6_0 & io_write_0_data_cf_loadWaitStrict | wenVec_6_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_6_cf_loadWaitBit = wenVec_6_0 & io_write_0_data_cf_loadWaitBit | wenVec_6_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2145 = wenVec_6_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2146 = wenVec_6_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_6_cf_waitForRobIdx_value = _wdata_T_2145 | _wdata_T_2146; // @[Mux.scala 27:73]
  wire  wdata_6_cf_waitForRobIdx_flag = wenVec_6_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_6_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_6_cf_storeSetHit = wenVec_6_0 & io_write_0_data_cf_storeSetHit | wenVec_6_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_6_cf_pred_taken = wenVec_6_0 & io_write_0_data_cf_pred_taken | wenVec_6_1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_6_cf_pd_isRet = wenVec_6_0 & io_write_0_data_cf_pd_isRet | wenVec_6_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_6_cf_pd_isCall = wenVec_6_0 & io_write_0_data_cf_pd_isCall | wenVec_6_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_2166 = wenVec_6_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_2167 = wenVec_6_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_6_cf_pd_brType = _wdata_T_2166 | _wdata_T_2167; // @[Mux.scala 27:73]
  wire  wdata_6_cf_pd_isRVC = wenVec_6_0 & io_write_0_data_cf_pd_isRVC | wenVec_6_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_6_cf_trigger_backendEn_0 = wenVec_6_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_6_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_6_cf_trigger_backendEn_1 = wenVec_6_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_6_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_2259 = wenVec_6_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_2260 = wenVec_6_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_6_cf_foldpc = _wdata_T_2259 | _wdata_T_2260; // @[Mux.scala 27:73]
  wire  wenVec_7_0 = io_write_0_enable & io_write_0_addr[7]; // @[PayloadArray.scala 55:53]
  wire  wenVec_7_1 = io_write_1_enable & io_write_1_addr[7]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_7 = {wenVec_7_1,wenVec_7_0}; // @[PayloadArray.scala 56:22]
  wire  wen_7 = |_wen_T_7; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_2301 = wenVec_7_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2302 = wenVec_7_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_7_sqIdx_value = _wdata_T_2301 | _wdata_T_2302; // @[Mux.scala 27:73]
  wire  wdata_7_sqIdx_flag = wenVec_7_0 & io_write_0_data_sqIdx_flag | wenVec_7_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2307 = wenVec_7_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2308 = wenVec_7_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_7_lqIdx_value = _wdata_T_2307 | _wdata_T_2308; // @[Mux.scala 27:73]
  wire  wdata_7_lqIdx_flag = wenVec_7_0 & io_write_0_data_lqIdx_flag | wenVec_7_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2313 = wenVec_7_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2314 = wenVec_7_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_7_robIdx_value = _wdata_T_2313 | _wdata_T_2314; // @[Mux.scala 27:73]
  wire  wdata_7_robIdx_flag = wenVec_7_0 & io_write_0_data_robIdx_flag | wenVec_7_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_2322 = wenVec_7_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_2323 = wenVec_7_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_7_pdest = _wdata_T_2322 | _wdata_T_2323; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_2397 = wenVec_7_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_2398 = wenVec_7_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_7_ctrl_imm = _wdata_T_2397 | _wdata_T_2398; // @[Mux.scala 27:73]
  wire  wdata_7_ctrl_fpWen = wenVec_7_0 & io_write_0_data_ctrl_fpWen | wenVec_7_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_7_ctrl_rfWen = wenVec_7_0 & io_write_0_data_ctrl_rfWen | wenVec_7_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_2421 = wenVec_7_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_2422 = wenVec_7_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_7_ctrl_fuOpType = _wdata_T_2421 | _wdata_T_2422; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2424 = wenVec_7_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2425 = wenVec_7_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_7_ctrl_fuType = _wdata_T_2424 | _wdata_T_2425; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2451 = wenVec_7_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2452 = wenVec_7_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_7_cf_ftqOffset = _wdata_T_2451 | _wdata_T_2452; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2454 = wenVec_7_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2455 = wenVec_7_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_7_cf_ftqPtr_value = _wdata_T_2454 | _wdata_T_2455; // @[Mux.scala 27:73]
  wire  wdata_7_cf_ftqPtr_flag = wenVec_7_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_7_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2460 = wenVec_7_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2461 = wenVec_7_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_7_cf_ssid = _wdata_T_2460 | _wdata_T_2461; // @[Mux.scala 27:73]
  wire  wdata_7_cf_loadWaitStrict = wenVec_7_0 & io_write_0_data_cf_loadWaitStrict | wenVec_7_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_7_cf_loadWaitBit = wenVec_7_0 & io_write_0_data_cf_loadWaitBit | wenVec_7_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2469 = wenVec_7_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2470 = wenVec_7_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_7_cf_waitForRobIdx_value = _wdata_T_2469 | _wdata_T_2470; // @[Mux.scala 27:73]
  wire  wdata_7_cf_waitForRobIdx_flag = wenVec_7_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_7_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_7_cf_storeSetHit = wenVec_7_0 & io_write_0_data_cf_storeSetHit | wenVec_7_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_7_cf_pred_taken = wenVec_7_0 & io_write_0_data_cf_pred_taken | wenVec_7_1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_7_cf_pd_isRet = wenVec_7_0 & io_write_0_data_cf_pd_isRet | wenVec_7_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_7_cf_pd_isCall = wenVec_7_0 & io_write_0_data_cf_pd_isCall | wenVec_7_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_2490 = wenVec_7_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_2491 = wenVec_7_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_7_cf_pd_brType = _wdata_T_2490 | _wdata_T_2491; // @[Mux.scala 27:73]
  wire  wdata_7_cf_pd_isRVC = wenVec_7_0 & io_write_0_data_cf_pd_isRVC | wenVec_7_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_7_cf_trigger_backendEn_0 = wenVec_7_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_7_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_7_cf_trigger_backendEn_1 = wenVec_7_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_7_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_2583 = wenVec_7_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_2584 = wenVec_7_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_7_cf_foldpc = _wdata_T_2583 | _wdata_T_2584; // @[Mux.scala 27:73]
  wire  wenVec_8_0 = io_write_0_enable & io_write_0_addr[8]; // @[PayloadArray.scala 55:53]
  wire  wenVec_8_1 = io_write_1_enable & io_write_1_addr[8]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_8 = {wenVec_8_1,wenVec_8_0}; // @[PayloadArray.scala 56:22]
  wire  wen_8 = |_wen_T_8; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_2625 = wenVec_8_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2626 = wenVec_8_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_8_sqIdx_value = _wdata_T_2625 | _wdata_T_2626; // @[Mux.scala 27:73]
  wire  wdata_8_sqIdx_flag = wenVec_8_0 & io_write_0_data_sqIdx_flag | wenVec_8_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2631 = wenVec_8_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2632 = wenVec_8_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_8_lqIdx_value = _wdata_T_2631 | _wdata_T_2632; // @[Mux.scala 27:73]
  wire  wdata_8_lqIdx_flag = wenVec_8_0 & io_write_0_data_lqIdx_flag | wenVec_8_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2637 = wenVec_8_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2638 = wenVec_8_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_8_robIdx_value = _wdata_T_2637 | _wdata_T_2638; // @[Mux.scala 27:73]
  wire  wdata_8_robIdx_flag = wenVec_8_0 & io_write_0_data_robIdx_flag | wenVec_8_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_2646 = wenVec_8_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_2647 = wenVec_8_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_8_pdest = _wdata_T_2646 | _wdata_T_2647; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_2721 = wenVec_8_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_2722 = wenVec_8_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_8_ctrl_imm = _wdata_T_2721 | _wdata_T_2722; // @[Mux.scala 27:73]
  wire  wdata_8_ctrl_fpWen = wenVec_8_0 & io_write_0_data_ctrl_fpWen | wenVec_8_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_8_ctrl_rfWen = wenVec_8_0 & io_write_0_data_ctrl_rfWen | wenVec_8_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_2745 = wenVec_8_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_2746 = wenVec_8_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_8_ctrl_fuOpType = _wdata_T_2745 | _wdata_T_2746; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2748 = wenVec_8_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2749 = wenVec_8_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_8_ctrl_fuType = _wdata_T_2748 | _wdata_T_2749; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2775 = wenVec_8_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2776 = wenVec_8_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_8_cf_ftqOffset = _wdata_T_2775 | _wdata_T_2776; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2778 = wenVec_8_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_2779 = wenVec_8_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_8_cf_ftqPtr_value = _wdata_T_2778 | _wdata_T_2779; // @[Mux.scala 27:73]
  wire  wdata_8_cf_ftqPtr_flag = wenVec_8_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_8_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2784 = wenVec_8_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2785 = wenVec_8_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_8_cf_ssid = _wdata_T_2784 | _wdata_T_2785; // @[Mux.scala 27:73]
  wire  wdata_8_cf_loadWaitStrict = wenVec_8_0 & io_write_0_data_cf_loadWaitStrict | wenVec_8_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_8_cf_loadWaitBit = wenVec_8_0 & io_write_0_data_cf_loadWaitBit | wenVec_8_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2793 = wenVec_8_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2794 = wenVec_8_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_8_cf_waitForRobIdx_value = _wdata_T_2793 | _wdata_T_2794; // @[Mux.scala 27:73]
  wire  wdata_8_cf_waitForRobIdx_flag = wenVec_8_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_8_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_8_cf_storeSetHit = wenVec_8_0 & io_write_0_data_cf_storeSetHit | wenVec_8_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_8_cf_pred_taken = wenVec_8_0 & io_write_0_data_cf_pred_taken | wenVec_8_1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_8_cf_pd_isRet = wenVec_8_0 & io_write_0_data_cf_pd_isRet | wenVec_8_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_8_cf_pd_isCall = wenVec_8_0 & io_write_0_data_cf_pd_isCall | wenVec_8_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_2814 = wenVec_8_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_2815 = wenVec_8_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_8_cf_pd_brType = _wdata_T_2814 | _wdata_T_2815; // @[Mux.scala 27:73]
  wire  wdata_8_cf_pd_isRVC = wenVec_8_0 & io_write_0_data_cf_pd_isRVC | wenVec_8_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_8_cf_trigger_backendEn_0 = wenVec_8_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_8_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_8_cf_trigger_backendEn_1 = wenVec_8_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_8_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_2907 = wenVec_8_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_2908 = wenVec_8_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_8_cf_foldpc = _wdata_T_2907 | _wdata_T_2908; // @[Mux.scala 27:73]
  wire  wenVec_9_0 = io_write_0_enable & io_write_0_addr[9]; // @[PayloadArray.scala 55:53]
  wire  wenVec_9_1 = io_write_1_enable & io_write_1_addr[9]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_9 = {wenVec_9_1,wenVec_9_0}; // @[PayloadArray.scala 56:22]
  wire  wen_9 = |_wen_T_9; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_2949 = wenVec_9_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2950 = wenVec_9_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_9_sqIdx_value = _wdata_T_2949 | _wdata_T_2950; // @[Mux.scala 27:73]
  wire  wdata_9_sqIdx_flag = wenVec_9_0 & io_write_0_data_sqIdx_flag | wenVec_9_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2955 = wenVec_9_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_2956 = wenVec_9_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_9_lqIdx_value = _wdata_T_2955 | _wdata_T_2956; // @[Mux.scala 27:73]
  wire  wdata_9_lqIdx_flag = wenVec_9_0 & io_write_0_data_lqIdx_flag | wenVec_9_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2961 = wenVec_9_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_2962 = wenVec_9_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_9_robIdx_value = _wdata_T_2961 | _wdata_T_2962; // @[Mux.scala 27:73]
  wire  wdata_9_robIdx_flag = wenVec_9_0 & io_write_0_data_robIdx_flag | wenVec_9_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_2970 = wenVec_9_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_2971 = wenVec_9_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_9_pdest = _wdata_T_2970 | _wdata_T_2971; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_3045 = wenVec_9_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_3046 = wenVec_9_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_9_ctrl_imm = _wdata_T_3045 | _wdata_T_3046; // @[Mux.scala 27:73]
  wire  wdata_9_ctrl_fpWen = wenVec_9_0 & io_write_0_data_ctrl_fpWen | wenVec_9_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_9_ctrl_rfWen = wenVec_9_0 & io_write_0_data_ctrl_rfWen | wenVec_9_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_3069 = wenVec_9_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_3070 = wenVec_9_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_9_ctrl_fuOpType = _wdata_T_3069 | _wdata_T_3070; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3072 = wenVec_9_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3073 = wenVec_9_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_9_ctrl_fuType = _wdata_T_3072 | _wdata_T_3073; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3099 = wenVec_9_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3100 = wenVec_9_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_9_cf_ftqOffset = _wdata_T_3099 | _wdata_T_3100; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3102 = wenVec_9_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3103 = wenVec_9_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_9_cf_ftqPtr_value = _wdata_T_3102 | _wdata_T_3103; // @[Mux.scala 27:73]
  wire  wdata_9_cf_ftqPtr_flag = wenVec_9_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_9_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3108 = wenVec_9_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3109 = wenVec_9_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_9_cf_ssid = _wdata_T_3108 | _wdata_T_3109; // @[Mux.scala 27:73]
  wire  wdata_9_cf_loadWaitStrict = wenVec_9_0 & io_write_0_data_cf_loadWaitStrict | wenVec_9_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_9_cf_loadWaitBit = wenVec_9_0 & io_write_0_data_cf_loadWaitBit | wenVec_9_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3117 = wenVec_9_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3118 = wenVec_9_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_9_cf_waitForRobIdx_value = _wdata_T_3117 | _wdata_T_3118; // @[Mux.scala 27:73]
  wire  wdata_9_cf_waitForRobIdx_flag = wenVec_9_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_9_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_9_cf_storeSetHit = wenVec_9_0 & io_write_0_data_cf_storeSetHit | wenVec_9_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_9_cf_pred_taken = wenVec_9_0 & io_write_0_data_cf_pred_taken | wenVec_9_1 & io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_9_cf_pd_isRet = wenVec_9_0 & io_write_0_data_cf_pd_isRet | wenVec_9_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_9_cf_pd_isCall = wenVec_9_0 & io_write_0_data_cf_pd_isCall | wenVec_9_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_3138 = wenVec_9_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_3139 = wenVec_9_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_9_cf_pd_brType = _wdata_T_3138 | _wdata_T_3139; // @[Mux.scala 27:73]
  wire  wdata_9_cf_pd_isRVC = wenVec_9_0 & io_write_0_data_cf_pd_isRVC | wenVec_9_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_9_cf_trigger_backendEn_0 = wenVec_9_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_9_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_9_cf_trigger_backendEn_1 = wenVec_9_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_9_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_3231 = wenVec_9_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_3232 = wenVec_9_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_9_cf_foldpc = _wdata_T_3231 | _wdata_T_3232; // @[Mux.scala 27:73]
  wire  wenVec_10_0 = io_write_0_enable & io_write_0_addr[10]; // @[PayloadArray.scala 55:53]
  wire  wenVec_10_1 = io_write_1_enable & io_write_1_addr[10]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_10 = {wenVec_10_1,wenVec_10_0}; // @[PayloadArray.scala 56:22]
  wire  wen_10 = |_wen_T_10; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_3273 = wenVec_10_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3274 = wenVec_10_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_10_sqIdx_value = _wdata_T_3273 | _wdata_T_3274; // @[Mux.scala 27:73]
  wire  wdata_10_sqIdx_flag = wenVec_10_0 & io_write_0_data_sqIdx_flag | wenVec_10_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3279 = wenVec_10_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3280 = wenVec_10_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_10_lqIdx_value = _wdata_T_3279 | _wdata_T_3280; // @[Mux.scala 27:73]
  wire  wdata_10_lqIdx_flag = wenVec_10_0 & io_write_0_data_lqIdx_flag | wenVec_10_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3285 = wenVec_10_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3286 = wenVec_10_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_10_robIdx_value = _wdata_T_3285 | _wdata_T_3286; // @[Mux.scala 27:73]
  wire  wdata_10_robIdx_flag = wenVec_10_0 & io_write_0_data_robIdx_flag | wenVec_10_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_3294 = wenVec_10_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_3295 = wenVec_10_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_10_pdest = _wdata_T_3294 | _wdata_T_3295; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_3369 = wenVec_10_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_3370 = wenVec_10_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_10_ctrl_imm = _wdata_T_3369 | _wdata_T_3370; // @[Mux.scala 27:73]
  wire  wdata_10_ctrl_fpWen = wenVec_10_0 & io_write_0_data_ctrl_fpWen | wenVec_10_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_10_ctrl_rfWen = wenVec_10_0 & io_write_0_data_ctrl_rfWen | wenVec_10_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_3393 = wenVec_10_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_3394 = wenVec_10_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_10_ctrl_fuOpType = _wdata_T_3393 | _wdata_T_3394; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3396 = wenVec_10_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3397 = wenVec_10_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_10_ctrl_fuType = _wdata_T_3396 | _wdata_T_3397; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3423 = wenVec_10_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3424 = wenVec_10_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_10_cf_ftqOffset = _wdata_T_3423 | _wdata_T_3424; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3426 = wenVec_10_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3427 = wenVec_10_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_10_cf_ftqPtr_value = _wdata_T_3426 | _wdata_T_3427; // @[Mux.scala 27:73]
  wire  wdata_10_cf_ftqPtr_flag = wenVec_10_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_10_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3432 = wenVec_10_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3433 = wenVec_10_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_10_cf_ssid = _wdata_T_3432 | _wdata_T_3433; // @[Mux.scala 27:73]
  wire  wdata_10_cf_loadWaitStrict = wenVec_10_0 & io_write_0_data_cf_loadWaitStrict | wenVec_10_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_10_cf_loadWaitBit = wenVec_10_0 & io_write_0_data_cf_loadWaitBit | wenVec_10_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3441 = wenVec_10_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3442 = wenVec_10_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_10_cf_waitForRobIdx_value = _wdata_T_3441 | _wdata_T_3442; // @[Mux.scala 27:73]
  wire  wdata_10_cf_waitForRobIdx_flag = wenVec_10_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_10_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_10_cf_storeSetHit = wenVec_10_0 & io_write_0_data_cf_storeSetHit | wenVec_10_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_10_cf_pred_taken = wenVec_10_0 & io_write_0_data_cf_pred_taken | wenVec_10_1 &
    io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_10_cf_pd_isRet = wenVec_10_0 & io_write_0_data_cf_pd_isRet | wenVec_10_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_10_cf_pd_isCall = wenVec_10_0 & io_write_0_data_cf_pd_isCall | wenVec_10_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_3462 = wenVec_10_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_3463 = wenVec_10_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_10_cf_pd_brType = _wdata_T_3462 | _wdata_T_3463; // @[Mux.scala 27:73]
  wire  wdata_10_cf_pd_isRVC = wenVec_10_0 & io_write_0_data_cf_pd_isRVC | wenVec_10_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_10_cf_trigger_backendEn_0 = wenVec_10_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_10_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_10_cf_trigger_backendEn_1 = wenVec_10_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_10_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_3555 = wenVec_10_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_3556 = wenVec_10_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_10_cf_foldpc = _wdata_T_3555 | _wdata_T_3556; // @[Mux.scala 27:73]
  wire  wenVec_11_0 = io_write_0_enable & io_write_0_addr[11]; // @[PayloadArray.scala 55:53]
  wire  wenVec_11_1 = io_write_1_enable & io_write_1_addr[11]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_11 = {wenVec_11_1,wenVec_11_0}; // @[PayloadArray.scala 56:22]
  wire  wen_11 = |_wen_T_11; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_3597 = wenVec_11_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3598 = wenVec_11_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_11_sqIdx_value = _wdata_T_3597 | _wdata_T_3598; // @[Mux.scala 27:73]
  wire  wdata_11_sqIdx_flag = wenVec_11_0 & io_write_0_data_sqIdx_flag | wenVec_11_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3603 = wenVec_11_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3604 = wenVec_11_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_11_lqIdx_value = _wdata_T_3603 | _wdata_T_3604; // @[Mux.scala 27:73]
  wire  wdata_11_lqIdx_flag = wenVec_11_0 & io_write_0_data_lqIdx_flag | wenVec_11_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3609 = wenVec_11_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3610 = wenVec_11_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_11_robIdx_value = _wdata_T_3609 | _wdata_T_3610; // @[Mux.scala 27:73]
  wire  wdata_11_robIdx_flag = wenVec_11_0 & io_write_0_data_robIdx_flag | wenVec_11_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_3618 = wenVec_11_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_3619 = wenVec_11_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_11_pdest = _wdata_T_3618 | _wdata_T_3619; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_3693 = wenVec_11_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_3694 = wenVec_11_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_11_ctrl_imm = _wdata_T_3693 | _wdata_T_3694; // @[Mux.scala 27:73]
  wire  wdata_11_ctrl_fpWen = wenVec_11_0 & io_write_0_data_ctrl_fpWen | wenVec_11_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_11_ctrl_rfWen = wenVec_11_0 & io_write_0_data_ctrl_rfWen | wenVec_11_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_3717 = wenVec_11_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_3718 = wenVec_11_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_11_ctrl_fuOpType = _wdata_T_3717 | _wdata_T_3718; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3720 = wenVec_11_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3721 = wenVec_11_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_11_ctrl_fuType = _wdata_T_3720 | _wdata_T_3721; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3747 = wenVec_11_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3748 = wenVec_11_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_11_cf_ftqOffset = _wdata_T_3747 | _wdata_T_3748; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3750 = wenVec_11_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_3751 = wenVec_11_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_11_cf_ftqPtr_value = _wdata_T_3750 | _wdata_T_3751; // @[Mux.scala 27:73]
  wire  wdata_11_cf_ftqPtr_flag = wenVec_11_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_11_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3756 = wenVec_11_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3757 = wenVec_11_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_11_cf_ssid = _wdata_T_3756 | _wdata_T_3757; // @[Mux.scala 27:73]
  wire  wdata_11_cf_loadWaitStrict = wenVec_11_0 & io_write_0_data_cf_loadWaitStrict | wenVec_11_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_11_cf_loadWaitBit = wenVec_11_0 & io_write_0_data_cf_loadWaitBit | wenVec_11_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3765 = wenVec_11_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3766 = wenVec_11_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_11_cf_waitForRobIdx_value = _wdata_T_3765 | _wdata_T_3766; // @[Mux.scala 27:73]
  wire  wdata_11_cf_waitForRobIdx_flag = wenVec_11_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_11_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_11_cf_storeSetHit = wenVec_11_0 & io_write_0_data_cf_storeSetHit | wenVec_11_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_11_cf_pred_taken = wenVec_11_0 & io_write_0_data_cf_pred_taken | wenVec_11_1 &
    io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_11_cf_pd_isRet = wenVec_11_0 & io_write_0_data_cf_pd_isRet | wenVec_11_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_11_cf_pd_isCall = wenVec_11_0 & io_write_0_data_cf_pd_isCall | wenVec_11_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_3786 = wenVec_11_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_3787 = wenVec_11_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_11_cf_pd_brType = _wdata_T_3786 | _wdata_T_3787; // @[Mux.scala 27:73]
  wire  wdata_11_cf_pd_isRVC = wenVec_11_0 & io_write_0_data_cf_pd_isRVC | wenVec_11_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_11_cf_trigger_backendEn_0 = wenVec_11_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_11_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_11_cf_trigger_backendEn_1 = wenVec_11_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_11_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_3879 = wenVec_11_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_3880 = wenVec_11_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_11_cf_foldpc = _wdata_T_3879 | _wdata_T_3880; // @[Mux.scala 27:73]
  wire  wenVec_12_0 = io_write_0_enable & io_write_0_addr[12]; // @[PayloadArray.scala 55:53]
  wire  wenVec_12_1 = io_write_1_enable & io_write_1_addr[12]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_12 = {wenVec_12_1,wenVec_12_0}; // @[PayloadArray.scala 56:22]
  wire  wen_12 = |_wen_T_12; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_3921 = wenVec_12_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3922 = wenVec_12_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_12_sqIdx_value = _wdata_T_3921 | _wdata_T_3922; // @[Mux.scala 27:73]
  wire  wdata_12_sqIdx_flag = wenVec_12_0 & io_write_0_data_sqIdx_flag | wenVec_12_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3927 = wenVec_12_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_3928 = wenVec_12_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_12_lqIdx_value = _wdata_T_3927 | _wdata_T_3928; // @[Mux.scala 27:73]
  wire  wdata_12_lqIdx_flag = wenVec_12_0 & io_write_0_data_lqIdx_flag | wenVec_12_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3933 = wenVec_12_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_3934 = wenVec_12_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_12_robIdx_value = _wdata_T_3933 | _wdata_T_3934; // @[Mux.scala 27:73]
  wire  wdata_12_robIdx_flag = wenVec_12_0 & io_write_0_data_robIdx_flag | wenVec_12_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_3942 = wenVec_12_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_3943 = wenVec_12_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_12_pdest = _wdata_T_3942 | _wdata_T_3943; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_4017 = wenVec_12_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_4018 = wenVec_12_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_12_ctrl_imm = _wdata_T_4017 | _wdata_T_4018; // @[Mux.scala 27:73]
  wire  wdata_12_ctrl_fpWen = wenVec_12_0 & io_write_0_data_ctrl_fpWen | wenVec_12_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_12_ctrl_rfWen = wenVec_12_0 & io_write_0_data_ctrl_rfWen | wenVec_12_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_4041 = wenVec_12_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_4042 = wenVec_12_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_12_ctrl_fuOpType = _wdata_T_4041 | _wdata_T_4042; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4044 = wenVec_12_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4045 = wenVec_12_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_12_ctrl_fuType = _wdata_T_4044 | _wdata_T_4045; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4071 = wenVec_12_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4072 = wenVec_12_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_12_cf_ftqOffset = _wdata_T_4071 | _wdata_T_4072; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4074 = wenVec_12_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4075 = wenVec_12_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_12_cf_ftqPtr_value = _wdata_T_4074 | _wdata_T_4075; // @[Mux.scala 27:73]
  wire  wdata_12_cf_ftqPtr_flag = wenVec_12_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_12_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4080 = wenVec_12_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4081 = wenVec_12_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_12_cf_ssid = _wdata_T_4080 | _wdata_T_4081; // @[Mux.scala 27:73]
  wire  wdata_12_cf_loadWaitStrict = wenVec_12_0 & io_write_0_data_cf_loadWaitStrict | wenVec_12_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_12_cf_loadWaitBit = wenVec_12_0 & io_write_0_data_cf_loadWaitBit | wenVec_12_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4089 = wenVec_12_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4090 = wenVec_12_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_12_cf_waitForRobIdx_value = _wdata_T_4089 | _wdata_T_4090; // @[Mux.scala 27:73]
  wire  wdata_12_cf_waitForRobIdx_flag = wenVec_12_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_12_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_12_cf_storeSetHit = wenVec_12_0 & io_write_0_data_cf_storeSetHit | wenVec_12_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_12_cf_pred_taken = wenVec_12_0 & io_write_0_data_cf_pred_taken | wenVec_12_1 &
    io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_12_cf_pd_isRet = wenVec_12_0 & io_write_0_data_cf_pd_isRet | wenVec_12_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_12_cf_pd_isCall = wenVec_12_0 & io_write_0_data_cf_pd_isCall | wenVec_12_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_4110 = wenVec_12_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_4111 = wenVec_12_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_12_cf_pd_brType = _wdata_T_4110 | _wdata_T_4111; // @[Mux.scala 27:73]
  wire  wdata_12_cf_pd_isRVC = wenVec_12_0 & io_write_0_data_cf_pd_isRVC | wenVec_12_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_12_cf_trigger_backendEn_0 = wenVec_12_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_12_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_12_cf_trigger_backendEn_1 = wenVec_12_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_12_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_4203 = wenVec_12_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_4204 = wenVec_12_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_12_cf_foldpc = _wdata_T_4203 | _wdata_T_4204; // @[Mux.scala 27:73]
  wire  wenVec_13_0 = io_write_0_enable & io_write_0_addr[13]; // @[PayloadArray.scala 55:53]
  wire  wenVec_13_1 = io_write_1_enable & io_write_1_addr[13]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_13 = {wenVec_13_1,wenVec_13_0}; // @[PayloadArray.scala 56:22]
  wire  wen_13 = |_wen_T_13; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_4245 = wenVec_13_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4246 = wenVec_13_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_13_sqIdx_value = _wdata_T_4245 | _wdata_T_4246; // @[Mux.scala 27:73]
  wire  wdata_13_sqIdx_flag = wenVec_13_0 & io_write_0_data_sqIdx_flag | wenVec_13_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4251 = wenVec_13_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4252 = wenVec_13_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_13_lqIdx_value = _wdata_T_4251 | _wdata_T_4252; // @[Mux.scala 27:73]
  wire  wdata_13_lqIdx_flag = wenVec_13_0 & io_write_0_data_lqIdx_flag | wenVec_13_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4257 = wenVec_13_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4258 = wenVec_13_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_13_robIdx_value = _wdata_T_4257 | _wdata_T_4258; // @[Mux.scala 27:73]
  wire  wdata_13_robIdx_flag = wenVec_13_0 & io_write_0_data_robIdx_flag | wenVec_13_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_4266 = wenVec_13_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_4267 = wenVec_13_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_13_pdest = _wdata_T_4266 | _wdata_T_4267; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_4341 = wenVec_13_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_4342 = wenVec_13_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_13_ctrl_imm = _wdata_T_4341 | _wdata_T_4342; // @[Mux.scala 27:73]
  wire  wdata_13_ctrl_fpWen = wenVec_13_0 & io_write_0_data_ctrl_fpWen | wenVec_13_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_13_ctrl_rfWen = wenVec_13_0 & io_write_0_data_ctrl_rfWen | wenVec_13_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_4365 = wenVec_13_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_4366 = wenVec_13_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_13_ctrl_fuOpType = _wdata_T_4365 | _wdata_T_4366; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4368 = wenVec_13_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4369 = wenVec_13_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_13_ctrl_fuType = _wdata_T_4368 | _wdata_T_4369; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4395 = wenVec_13_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4396 = wenVec_13_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_13_cf_ftqOffset = _wdata_T_4395 | _wdata_T_4396; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4398 = wenVec_13_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4399 = wenVec_13_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_13_cf_ftqPtr_value = _wdata_T_4398 | _wdata_T_4399; // @[Mux.scala 27:73]
  wire  wdata_13_cf_ftqPtr_flag = wenVec_13_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_13_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4404 = wenVec_13_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4405 = wenVec_13_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_13_cf_ssid = _wdata_T_4404 | _wdata_T_4405; // @[Mux.scala 27:73]
  wire  wdata_13_cf_loadWaitStrict = wenVec_13_0 & io_write_0_data_cf_loadWaitStrict | wenVec_13_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_13_cf_loadWaitBit = wenVec_13_0 & io_write_0_data_cf_loadWaitBit | wenVec_13_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4413 = wenVec_13_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4414 = wenVec_13_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_13_cf_waitForRobIdx_value = _wdata_T_4413 | _wdata_T_4414; // @[Mux.scala 27:73]
  wire  wdata_13_cf_waitForRobIdx_flag = wenVec_13_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_13_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_13_cf_storeSetHit = wenVec_13_0 & io_write_0_data_cf_storeSetHit | wenVec_13_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_13_cf_pred_taken = wenVec_13_0 & io_write_0_data_cf_pred_taken | wenVec_13_1 &
    io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_13_cf_pd_isRet = wenVec_13_0 & io_write_0_data_cf_pd_isRet | wenVec_13_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_13_cf_pd_isCall = wenVec_13_0 & io_write_0_data_cf_pd_isCall | wenVec_13_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_4434 = wenVec_13_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_4435 = wenVec_13_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_13_cf_pd_brType = _wdata_T_4434 | _wdata_T_4435; // @[Mux.scala 27:73]
  wire  wdata_13_cf_pd_isRVC = wenVec_13_0 & io_write_0_data_cf_pd_isRVC | wenVec_13_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_13_cf_trigger_backendEn_0 = wenVec_13_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_13_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_13_cf_trigger_backendEn_1 = wenVec_13_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_13_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_4527 = wenVec_13_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_4528 = wenVec_13_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_13_cf_foldpc = _wdata_T_4527 | _wdata_T_4528; // @[Mux.scala 27:73]
  wire  wenVec_14_0 = io_write_0_enable & io_write_0_addr[14]; // @[PayloadArray.scala 55:53]
  wire  wenVec_14_1 = io_write_1_enable & io_write_1_addr[14]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_14 = {wenVec_14_1,wenVec_14_0}; // @[PayloadArray.scala 56:22]
  wire  wen_14 = |_wen_T_14; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_4569 = wenVec_14_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4570 = wenVec_14_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_14_sqIdx_value = _wdata_T_4569 | _wdata_T_4570; // @[Mux.scala 27:73]
  wire  wdata_14_sqIdx_flag = wenVec_14_0 & io_write_0_data_sqIdx_flag | wenVec_14_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4575 = wenVec_14_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4576 = wenVec_14_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_14_lqIdx_value = _wdata_T_4575 | _wdata_T_4576; // @[Mux.scala 27:73]
  wire  wdata_14_lqIdx_flag = wenVec_14_0 & io_write_0_data_lqIdx_flag | wenVec_14_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4581 = wenVec_14_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4582 = wenVec_14_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_14_robIdx_value = _wdata_T_4581 | _wdata_T_4582; // @[Mux.scala 27:73]
  wire  wdata_14_robIdx_flag = wenVec_14_0 & io_write_0_data_robIdx_flag | wenVec_14_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_4590 = wenVec_14_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_4591 = wenVec_14_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_14_pdest = _wdata_T_4590 | _wdata_T_4591; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_4665 = wenVec_14_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_4666 = wenVec_14_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_14_ctrl_imm = _wdata_T_4665 | _wdata_T_4666; // @[Mux.scala 27:73]
  wire  wdata_14_ctrl_fpWen = wenVec_14_0 & io_write_0_data_ctrl_fpWen | wenVec_14_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_14_ctrl_rfWen = wenVec_14_0 & io_write_0_data_ctrl_rfWen | wenVec_14_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_4689 = wenVec_14_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_4690 = wenVec_14_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_14_ctrl_fuOpType = _wdata_T_4689 | _wdata_T_4690; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4692 = wenVec_14_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4693 = wenVec_14_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_14_ctrl_fuType = _wdata_T_4692 | _wdata_T_4693; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4719 = wenVec_14_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4720 = wenVec_14_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_14_cf_ftqOffset = _wdata_T_4719 | _wdata_T_4720; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4722 = wenVec_14_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_4723 = wenVec_14_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_14_cf_ftqPtr_value = _wdata_T_4722 | _wdata_T_4723; // @[Mux.scala 27:73]
  wire  wdata_14_cf_ftqPtr_flag = wenVec_14_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_14_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4728 = wenVec_14_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4729 = wenVec_14_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_14_cf_ssid = _wdata_T_4728 | _wdata_T_4729; // @[Mux.scala 27:73]
  wire  wdata_14_cf_loadWaitStrict = wenVec_14_0 & io_write_0_data_cf_loadWaitStrict | wenVec_14_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_14_cf_loadWaitBit = wenVec_14_0 & io_write_0_data_cf_loadWaitBit | wenVec_14_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4737 = wenVec_14_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4738 = wenVec_14_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_14_cf_waitForRobIdx_value = _wdata_T_4737 | _wdata_T_4738; // @[Mux.scala 27:73]
  wire  wdata_14_cf_waitForRobIdx_flag = wenVec_14_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_14_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_14_cf_storeSetHit = wenVec_14_0 & io_write_0_data_cf_storeSetHit | wenVec_14_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_14_cf_pred_taken = wenVec_14_0 & io_write_0_data_cf_pred_taken | wenVec_14_1 &
    io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_14_cf_pd_isRet = wenVec_14_0 & io_write_0_data_cf_pd_isRet | wenVec_14_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_14_cf_pd_isCall = wenVec_14_0 & io_write_0_data_cf_pd_isCall | wenVec_14_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_4758 = wenVec_14_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_4759 = wenVec_14_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_14_cf_pd_brType = _wdata_T_4758 | _wdata_T_4759; // @[Mux.scala 27:73]
  wire  wdata_14_cf_pd_isRVC = wenVec_14_0 & io_write_0_data_cf_pd_isRVC | wenVec_14_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_14_cf_trigger_backendEn_0 = wenVec_14_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_14_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_14_cf_trigger_backendEn_1 = wenVec_14_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_14_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_4851 = wenVec_14_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_4852 = wenVec_14_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_14_cf_foldpc = _wdata_T_4851 | _wdata_T_4852; // @[Mux.scala 27:73]
  wire  wenVec_15_0 = io_write_0_enable & io_write_0_addr[15]; // @[PayloadArray.scala 55:53]
  wire  wenVec_15_1 = io_write_1_enable & io_write_1_addr[15]; // @[PayloadArray.scala 55:53]
  wire [1:0] _wen_T_15 = {wenVec_15_1,wenVec_15_0}; // @[PayloadArray.scala 56:22]
  wire  wen_15 = |_wen_T_15; // @[PayloadArray.scala 56:29]
  wire [3:0] _wdata_T_4893 = wenVec_15_0 ? io_write_0_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4894 = wenVec_15_1 ? io_write_1_data_sqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_15_sqIdx_value = _wdata_T_4893 | _wdata_T_4894; // @[Mux.scala 27:73]
  wire  wdata_15_sqIdx_flag = wenVec_15_0 & io_write_0_data_sqIdx_flag | wenVec_15_1 & io_write_1_data_sqIdx_flag; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4899 = wenVec_15_0 ? io_write_0_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_4900 = wenVec_15_1 ? io_write_1_data_lqIdx_value : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_15_lqIdx_value = _wdata_T_4899 | _wdata_T_4900; // @[Mux.scala 27:73]
  wire  wdata_15_lqIdx_flag = wenVec_15_0 & io_write_0_data_lqIdx_flag | wenVec_15_1 & io_write_1_data_lqIdx_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4905 = wenVec_15_0 ? io_write_0_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_4906 = wenVec_15_1 ? io_write_1_data_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_15_robIdx_value = _wdata_T_4905 | _wdata_T_4906; // @[Mux.scala 27:73]
  wire  wdata_15_robIdx_flag = wenVec_15_0 & io_write_0_data_robIdx_flag | wenVec_15_1 & io_write_1_data_robIdx_flag; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_4914 = wenVec_15_0 ? io_write_0_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _wdata_T_4915 = wenVec_15_1 ? io_write_1_data_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] wdata_15_pdest = _wdata_T_4914 | _wdata_T_4915; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_4989 = wenVec_15_0 ? io_write_0_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _wdata_T_4990 = wenVec_15_1 ? io_write_1_data_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] wdata_15_ctrl_imm = _wdata_T_4989 | _wdata_T_4990; // @[Mux.scala 27:73]
  wire  wdata_15_ctrl_fpWen = wenVec_15_0 & io_write_0_data_ctrl_fpWen | wenVec_15_1 & io_write_1_data_ctrl_fpWen; // @[Mux.scala 27:73]
  wire  wdata_15_ctrl_rfWen = wenVec_15_0 & io_write_0_data_ctrl_rfWen | wenVec_15_1 & io_write_1_data_ctrl_rfWen; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_5013 = wenVec_15_0 ? io_write_0_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _wdata_T_5014 = wenVec_15_1 ? io_write_1_data_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] wdata_15_ctrl_fuOpType = _wdata_T_5013 | _wdata_T_5014; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_5016 = wenVec_15_0 ? io_write_0_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _wdata_T_5017 = wenVec_15_1 ? io_write_1_data_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] wdata_15_ctrl_fuType = _wdata_T_5016 | _wdata_T_5017; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_5043 = wenVec_15_0 ? io_write_0_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_5044 = wenVec_15_1 ? io_write_1_data_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_15_cf_ftqOffset = _wdata_T_5043 | _wdata_T_5044; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_5046 = wenVec_15_0 ? io_write_0_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _wdata_T_5047 = wenVec_15_1 ? io_write_1_data_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] wdata_15_cf_ftqPtr_value = _wdata_T_5046 | _wdata_T_5047; // @[Mux.scala 27:73]
  wire  wdata_15_cf_ftqPtr_flag = wenVec_15_0 & io_write_0_data_cf_ftqPtr_flag | wenVec_15_1 &
    io_write_1_data_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_5052 = wenVec_15_0 ? io_write_0_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_5053 = wenVec_15_1 ? io_write_1_data_cf_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_15_cf_ssid = _wdata_T_5052 | _wdata_T_5053; // @[Mux.scala 27:73]
  wire  wdata_15_cf_loadWaitStrict = wenVec_15_0 & io_write_0_data_cf_loadWaitStrict | wenVec_15_1 &
    io_write_1_data_cf_loadWaitStrict; // @[Mux.scala 27:73]
  wire  wdata_15_cf_loadWaitBit = wenVec_15_0 & io_write_0_data_cf_loadWaitBit | wenVec_15_1 &
    io_write_1_data_cf_loadWaitBit; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_5061 = wenVec_15_0 ? io_write_0_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _wdata_T_5062 = wenVec_15_1 ? io_write_1_data_cf_waitForRobIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] wdata_15_cf_waitForRobIdx_value = _wdata_T_5061 | _wdata_T_5062; // @[Mux.scala 27:73]
  wire  wdata_15_cf_waitForRobIdx_flag = wenVec_15_0 & io_write_0_data_cf_waitForRobIdx_flag | wenVec_15_1 &
    io_write_1_data_cf_waitForRobIdx_flag; // @[Mux.scala 27:73]
  wire  wdata_15_cf_storeSetHit = wenVec_15_0 & io_write_0_data_cf_storeSetHit | wenVec_15_1 &
    io_write_1_data_cf_storeSetHit; // @[Mux.scala 27:73]
  wire  wdata_15_cf_pred_taken = wenVec_15_0 & io_write_0_data_cf_pred_taken | wenVec_15_1 &
    io_write_1_data_cf_pred_taken; // @[Mux.scala 27:73]
  wire  wdata_15_cf_pd_isRet = wenVec_15_0 & io_write_0_data_cf_pd_isRet | wenVec_15_1 & io_write_1_data_cf_pd_isRet; // @[Mux.scala 27:73]
  wire  wdata_15_cf_pd_isCall = wenVec_15_0 & io_write_0_data_cf_pd_isCall | wenVec_15_1 & io_write_1_data_cf_pd_isCall; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_5082 = wenVec_15_0 ? io_write_0_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _wdata_T_5083 = wenVec_15_1 ? io_write_1_data_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] wdata_15_cf_pd_brType = _wdata_T_5082 | _wdata_T_5083; // @[Mux.scala 27:73]
  wire  wdata_15_cf_pd_isRVC = wenVec_15_0 & io_write_0_data_cf_pd_isRVC | wenVec_15_1 & io_write_1_data_cf_pd_isRVC; // @[Mux.scala 27:73]
  wire  wdata_15_cf_trigger_backendEn_0 = wenVec_15_0 & io_write_0_data_cf_trigger_backendEn_0 | wenVec_15_1 &
    io_write_1_data_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  wire  wdata_15_cf_trigger_backendEn_1 = wenVec_15_0 & io_write_0_data_cf_trigger_backendEn_1 | wenVec_15_1 &
    io_write_1_data_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_5175 = wenVec_15_0 ? io_write_0_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _wdata_T_5176 = wenVec_15_1 ? io_write_1_data_cf_foldpc : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] wdata_15_cf_foldpc = _wdata_T_5175 | _wdata_T_5176; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_foldpc = _io_read_0_data_T_3300 | _io_read_0_data_T_3286; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_trigger_backendEn_0 = io_read_0_addr[0] & payload_0_cf_trigger_backendEn_0 | io_read_0_addr[1
    ] & payload_1_cf_trigger_backendEn_0 | io_read_0_addr[2] & payload_2_cf_trigger_backendEn_0 | io_read_0_addr[3] &
    payload_3_cf_trigger_backendEn_0 | io_read_0_addr[4] & payload_4_cf_trigger_backendEn_0 | io_read_0_addr[5] &
    payload_5_cf_trigger_backendEn_0 | io_read_0_addr[6] & payload_6_cf_trigger_backendEn_0 | io_read_0_addr[7] &
    payload_7_cf_trigger_backendEn_0 | io_read_0_addr[8] & payload_8_cf_trigger_backendEn_0 | io_read_0_addr[9] &
    payload_9_cf_trigger_backendEn_0 | io_read_0_addr[10] & payload_10_cf_trigger_backendEn_0 | io_read_0_addr[11] &
    payload_11_cf_trigger_backendEn_0 | io_read_0_addr[12] & payload_12_cf_trigger_backendEn_0 | io_read_0_addr[13] &
    payload_13_cf_trigger_backendEn_0 | io_read_0_addr[14] & payload_14_cf_trigger_backendEn_0 | _io_read_0_data_T_2604; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_trigger_backendEn_1 = io_read_0_addr[0] & payload_0_cf_trigger_backendEn_1 | io_read_0_addr[1
    ] & payload_1_cf_trigger_backendEn_1 | io_read_0_addr[2] & payload_2_cf_trigger_backendEn_1 | io_read_0_addr[3] &
    payload_3_cf_trigger_backendEn_1 | io_read_0_addr[4] & payload_4_cf_trigger_backendEn_1 | io_read_0_addr[5] &
    payload_5_cf_trigger_backendEn_1 | io_read_0_addr[6] & payload_6_cf_trigger_backendEn_1 | io_read_0_addr[7] &
    payload_7_cf_trigger_backendEn_1 | io_read_0_addr[8] & payload_8_cf_trigger_backendEn_1 | io_read_0_addr[9] &
    payload_9_cf_trigger_backendEn_1 | io_read_0_addr[10] & payload_10_cf_trigger_backendEn_1 | io_read_0_addr[11] &
    payload_11_cf_trigger_backendEn_1 | io_read_0_addr[12] & payload_12_cf_trigger_backendEn_1 | io_read_0_addr[13] &
    payload_13_cf_trigger_backendEn_1 | io_read_0_addr[14] & payload_14_cf_trigger_backendEn_1 | _io_read_0_data_T_2635; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_pd_isRVC = io_read_0_addr[0] & payload_0_cf_pd_isRVC | io_read_0_addr[1] &
    payload_1_cf_pd_isRVC | io_read_0_addr[2] & payload_2_cf_pd_isRVC | io_read_0_addr[3] & payload_3_cf_pd_isRVC |
    io_read_0_addr[4] & payload_4_cf_pd_isRVC | io_read_0_addr[5] & payload_5_cf_pd_isRVC | io_read_0_addr[6] &
    payload_6_cf_pd_isRVC | io_read_0_addr[7] & payload_7_cf_pd_isRVC | io_read_0_addr[8] & payload_8_cf_pd_isRVC |
    io_read_0_addr[9] & payload_9_cf_pd_isRVC | io_read_0_addr[10] & payload_10_cf_pd_isRVC | io_read_0_addr[11] &
    payload_11_cf_pd_isRVC | io_read_0_addr[12] & payload_12_cf_pd_isRVC | io_read_0_addr[13] & payload_13_cf_pd_isRVC
     | io_read_0_addr[14] & payload_14_cf_pd_isRVC | _io_read_0_data_T_2356; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_pd_brType = _io_read_0_data_T_2339 | _io_read_0_data_T_2325; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_pd_isCall = io_read_0_addr[0] & payload_0_cf_pd_isCall | io_read_0_addr[1] &
    payload_1_cf_pd_isCall | io_read_0_addr[2] & payload_2_cf_pd_isCall | io_read_0_addr[3] & payload_3_cf_pd_isCall |
    io_read_0_addr[4] & payload_4_cf_pd_isCall | io_read_0_addr[5] & payload_5_cf_pd_isCall | io_read_0_addr[6] &
    payload_6_cf_pd_isCall | io_read_0_addr[7] & payload_7_cf_pd_isCall | io_read_0_addr[8] & payload_8_cf_pd_isCall |
    io_read_0_addr[9] & payload_9_cf_pd_isCall | io_read_0_addr[10] & payload_10_cf_pd_isCall | io_read_0_addr[11] &
    payload_11_cf_pd_isCall | io_read_0_addr[12] & payload_12_cf_pd_isCall | io_read_0_addr[13] &
    payload_13_cf_pd_isCall | io_read_0_addr[14] & payload_14_cf_pd_isCall | _io_read_0_data_T_2294; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_pd_isRet = io_read_0_addr[0] & payload_0_cf_pd_isRet | io_read_0_addr[1] &
    payload_1_cf_pd_isRet | io_read_0_addr[2] & payload_2_cf_pd_isRet | io_read_0_addr[3] & payload_3_cf_pd_isRet |
    io_read_0_addr[4] & payload_4_cf_pd_isRet | io_read_0_addr[5] & payload_5_cf_pd_isRet | io_read_0_addr[6] &
    payload_6_cf_pd_isRet | io_read_0_addr[7] & payload_7_cf_pd_isRet | io_read_0_addr[8] & payload_8_cf_pd_isRet |
    io_read_0_addr[9] & payload_9_cf_pd_isRet | io_read_0_addr[10] & payload_10_cf_pd_isRet | io_read_0_addr[11] &
    payload_11_cf_pd_isRet | io_read_0_addr[12] & payload_12_cf_pd_isRet | io_read_0_addr[13] & payload_13_cf_pd_isRet
     | io_read_0_addr[14] & payload_14_cf_pd_isRet | _io_read_0_data_T_2263; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_pred_taken = io_read_0_addr[0] & payload_0_cf_pred_taken | io_read_0_addr[1] &
    payload_1_cf_pred_taken | io_read_0_addr[2] & payload_2_cf_pred_taken | io_read_0_addr[3] & payload_3_cf_pred_taken
     | io_read_0_addr[4] & payload_4_cf_pred_taken | io_read_0_addr[5] & payload_5_cf_pred_taken | io_read_0_addr[6] &
    payload_6_cf_pred_taken | io_read_0_addr[7] & payload_7_cf_pred_taken | io_read_0_addr[8] & payload_8_cf_pred_taken
     | io_read_0_addr[9] & payload_9_cf_pred_taken | io_read_0_addr[10] & payload_10_cf_pred_taken | io_read_0_addr[11]
     & payload_11_cf_pred_taken | io_read_0_addr[12] & payload_12_cf_pred_taken | io_read_0_addr[13] &
    payload_13_cf_pred_taken | io_read_0_addr[14] & payload_14_cf_pred_taken | _io_read_0_data_T_2232; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_storeSetHit = io_read_0_addr[0] & payload_0_cf_storeSetHit | io_read_0_addr[1] &
    payload_1_cf_storeSetHit | io_read_0_addr[2] & payload_2_cf_storeSetHit | io_read_0_addr[3] &
    payload_3_cf_storeSetHit | io_read_0_addr[4] & payload_4_cf_storeSetHit | io_read_0_addr[5] &
    payload_5_cf_storeSetHit | io_read_0_addr[6] & payload_6_cf_storeSetHit | io_read_0_addr[7] &
    payload_7_cf_storeSetHit | io_read_0_addr[8] & payload_8_cf_storeSetHit | io_read_0_addr[9] &
    payload_9_cf_storeSetHit | io_read_0_addr[10] & payload_10_cf_storeSetHit | io_read_0_addr[11] &
    payload_11_cf_storeSetHit | io_read_0_addr[12] & payload_12_cf_storeSetHit | io_read_0_addr[13] &
    payload_13_cf_storeSetHit | io_read_0_addr[14] & payload_14_cf_storeSetHit | _io_read_0_data_T_2170; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_waitForRobIdx_flag = io_read_0_addr[0] & payload_0_cf_waitForRobIdx_flag | io_read_0_addr[1]
     & payload_1_cf_waitForRobIdx_flag | io_read_0_addr[2] & payload_2_cf_waitForRobIdx_flag | io_read_0_addr[3] &
    payload_3_cf_waitForRobIdx_flag | io_read_0_addr[4] & payload_4_cf_waitForRobIdx_flag | io_read_0_addr[5] &
    payload_5_cf_waitForRobIdx_flag | io_read_0_addr[6] & payload_6_cf_waitForRobIdx_flag | io_read_0_addr[7] &
    payload_7_cf_waitForRobIdx_flag | io_read_0_addr[8] & payload_8_cf_waitForRobIdx_flag | io_read_0_addr[9] &
    payload_9_cf_waitForRobIdx_flag | io_read_0_addr[10] & payload_10_cf_waitForRobIdx_flag | io_read_0_addr[11] &
    payload_11_cf_waitForRobIdx_flag | io_read_0_addr[12] & payload_12_cf_waitForRobIdx_flag | io_read_0_addr[13] &
    payload_13_cf_waitForRobIdx_flag | io_read_0_addr[14] & payload_14_cf_waitForRobIdx_flag | _io_read_0_data_T_2139; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_waitForRobIdx_value = _io_read_0_data_T_2122 | _io_read_0_data_T_2108; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_loadWaitBit = io_read_0_addr[0] & payload_0_cf_loadWaitBit | io_read_0_addr[1] &
    payload_1_cf_loadWaitBit | io_read_0_addr[2] & payload_2_cf_loadWaitBit | io_read_0_addr[3] &
    payload_3_cf_loadWaitBit | io_read_0_addr[4] & payload_4_cf_loadWaitBit | io_read_0_addr[5] &
    payload_5_cf_loadWaitBit | io_read_0_addr[6] & payload_6_cf_loadWaitBit | io_read_0_addr[7] &
    payload_7_cf_loadWaitBit | io_read_0_addr[8] & payload_8_cf_loadWaitBit | io_read_0_addr[9] &
    payload_9_cf_loadWaitBit | io_read_0_addr[10] & payload_10_cf_loadWaitBit | io_read_0_addr[11] &
    payload_11_cf_loadWaitBit | io_read_0_addr[12] & payload_12_cf_loadWaitBit | io_read_0_addr[13] &
    payload_13_cf_loadWaitBit | io_read_0_addr[14] & payload_14_cf_loadWaitBit | _io_read_0_data_T_2077; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_loadWaitStrict = io_read_0_addr[0] & payload_0_cf_loadWaitStrict | io_read_0_addr[1] &
    payload_1_cf_loadWaitStrict | io_read_0_addr[2] & payload_2_cf_loadWaitStrict | io_read_0_addr[3] &
    payload_3_cf_loadWaitStrict | io_read_0_addr[4] & payload_4_cf_loadWaitStrict | io_read_0_addr[5] &
    payload_5_cf_loadWaitStrict | io_read_0_addr[6] & payload_6_cf_loadWaitStrict | io_read_0_addr[7] &
    payload_7_cf_loadWaitStrict | io_read_0_addr[8] & payload_8_cf_loadWaitStrict | io_read_0_addr[9] &
    payload_9_cf_loadWaitStrict | io_read_0_addr[10] & payload_10_cf_loadWaitStrict | io_read_0_addr[11] &
    payload_11_cf_loadWaitStrict | io_read_0_addr[12] & payload_12_cf_loadWaitStrict | io_read_0_addr[13] &
    payload_13_cf_loadWaitStrict | io_read_0_addr[14] & payload_14_cf_loadWaitStrict | _io_read_0_data_T_2046; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_ssid = _io_read_0_data_T_2029 | _io_read_0_data_T_2015; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_ftqPtr_flag = io_read_0_addr[0] & payload_0_cf_ftqPtr_flag | io_read_0_addr[1] &
    payload_1_cf_ftqPtr_flag | io_read_0_addr[2] & payload_2_cf_ftqPtr_flag | io_read_0_addr[3] &
    payload_3_cf_ftqPtr_flag | io_read_0_addr[4] & payload_4_cf_ftqPtr_flag | io_read_0_addr[5] &
    payload_5_cf_ftqPtr_flag | io_read_0_addr[6] & payload_6_cf_ftqPtr_flag | io_read_0_addr[7] &
    payload_7_cf_ftqPtr_flag | io_read_0_addr[8] & payload_8_cf_ftqPtr_flag | io_read_0_addr[9] &
    payload_9_cf_ftqPtr_flag | io_read_0_addr[10] & payload_10_cf_ftqPtr_flag | io_read_0_addr[11] &
    payload_11_cf_ftqPtr_flag | io_read_0_addr[12] & payload_12_cf_ftqPtr_flag | io_read_0_addr[13] &
    payload_13_cf_ftqPtr_flag | io_read_0_addr[14] & payload_14_cf_ftqPtr_flag | _io_read_0_data_T_1984; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_ftqPtr_value = _io_read_0_data_T_1967 | _io_read_0_data_T_1953; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_ftqOffset = _io_read_0_data_T_1936 | _io_read_0_data_T_1922; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fuType = _io_read_0_data_T_1657 | _io_read_0_data_T_1643; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fuOpType = _io_read_0_data_T_1626 | _io_read_0_data_T_1612; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_rfWen = io_read_0_addr[0] & payload_0_ctrl_rfWen | io_read_0_addr[1] & payload_1_ctrl_rfWen
     | io_read_0_addr[2] & payload_2_ctrl_rfWen | io_read_0_addr[3] & payload_3_ctrl_rfWen | io_read_0_addr[4] &
    payload_4_ctrl_rfWen | io_read_0_addr[5] & payload_5_ctrl_rfWen | io_read_0_addr[6] & payload_6_ctrl_rfWen |
    io_read_0_addr[7] & payload_7_ctrl_rfWen | io_read_0_addr[8] & payload_8_ctrl_rfWen | io_read_0_addr[9] &
    payload_9_ctrl_rfWen | io_read_0_addr[10] & payload_10_ctrl_rfWen | io_read_0_addr[11] & payload_11_ctrl_rfWen |
    io_read_0_addr[12] & payload_12_ctrl_rfWen | io_read_0_addr[13] & payload_13_ctrl_rfWen | io_read_0_addr[14] &
    payload_14_ctrl_rfWen | _io_read_0_data_T_1581; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpWen = io_read_0_addr[0] & payload_0_ctrl_fpWen | io_read_0_addr[1] & payload_1_ctrl_fpWen
     | io_read_0_addr[2] & payload_2_ctrl_fpWen | io_read_0_addr[3] & payload_3_ctrl_fpWen | io_read_0_addr[4] &
    payload_4_ctrl_fpWen | io_read_0_addr[5] & payload_5_ctrl_fpWen | io_read_0_addr[6] & payload_6_ctrl_fpWen |
    io_read_0_addr[7] & payload_7_ctrl_fpWen | io_read_0_addr[8] & payload_8_ctrl_fpWen | io_read_0_addr[9] &
    payload_9_ctrl_fpWen | io_read_0_addr[10] & payload_10_ctrl_fpWen | io_read_0_addr[11] & payload_11_ctrl_fpWen |
    io_read_0_addr[12] & payload_12_ctrl_fpWen | io_read_0_addr[13] & payload_13_ctrl_fpWen | io_read_0_addr[14] &
    payload_14_ctrl_fpWen | _io_read_0_data_T_1550; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_imm = _io_read_0_data_T_1378 | _io_read_0_data_T_1364; // @[Mux.scala 27:73]
  assign io_read_0_data_pdest = _io_read_0_data_T_603 | _io_read_0_data_T_589; // @[Mux.scala 27:73]
  assign io_read_0_data_robIdx_flag = io_read_0_addr[0] & payload_0_robIdx_flag | io_read_0_addr[1] &
    payload_1_robIdx_flag | io_read_0_addr[2] & payload_2_robIdx_flag | io_read_0_addr[3] & payload_3_robIdx_flag |
    io_read_0_addr[4] & payload_4_robIdx_flag | io_read_0_addr[5] & payload_5_robIdx_flag | io_read_0_addr[6] &
    payload_6_robIdx_flag | io_read_0_addr[7] & payload_7_robIdx_flag | io_read_0_addr[8] & payload_8_robIdx_flag |
    io_read_0_addr[9] & payload_9_robIdx_flag | io_read_0_addr[10] & payload_10_robIdx_flag | io_read_0_addr[11] &
    payload_11_robIdx_flag | io_read_0_addr[12] & payload_12_robIdx_flag | io_read_0_addr[13] & payload_13_robIdx_flag
     | io_read_0_addr[14] & payload_14_robIdx_flag | _io_read_0_data_T_527; // @[Mux.scala 27:73]
  assign io_read_0_data_robIdx_value = _io_read_0_data_T_510 | _io_read_0_data_T_496; // @[Mux.scala 27:73]
  assign io_read_0_data_lqIdx_flag = io_read_0_addr[0] & payload_0_lqIdx_flag | io_read_0_addr[1] & payload_1_lqIdx_flag
     | io_read_0_addr[2] & payload_2_lqIdx_flag | io_read_0_addr[3] & payload_3_lqIdx_flag | io_read_0_addr[4] &
    payload_4_lqIdx_flag | io_read_0_addr[5] & payload_5_lqIdx_flag | io_read_0_addr[6] & payload_6_lqIdx_flag |
    io_read_0_addr[7] & payload_7_lqIdx_flag | io_read_0_addr[8] & payload_8_lqIdx_flag | io_read_0_addr[9] &
    payload_9_lqIdx_flag | io_read_0_addr[10] & payload_10_lqIdx_flag | io_read_0_addr[11] & payload_11_lqIdx_flag |
    io_read_0_addr[12] & payload_12_lqIdx_flag | io_read_0_addr[13] & payload_13_lqIdx_flag | io_read_0_addr[14] &
    payload_14_lqIdx_flag | _io_read_0_data_T_465; // @[Mux.scala 27:73]
  assign io_read_0_data_lqIdx_value = _io_read_0_data_T_448 | _io_read_0_data_T_434; // @[Mux.scala 27:73]
  assign io_read_0_data_sqIdx_flag = io_read_0_addr[0] & payload_0_sqIdx_flag | io_read_0_addr[1] & payload_1_sqIdx_flag
     | io_read_0_addr[2] & payload_2_sqIdx_flag | io_read_0_addr[3] & payload_3_sqIdx_flag | io_read_0_addr[4] &
    payload_4_sqIdx_flag | io_read_0_addr[5] & payload_5_sqIdx_flag | io_read_0_addr[6] & payload_6_sqIdx_flag |
    io_read_0_addr[7] & payload_7_sqIdx_flag | io_read_0_addr[8] & payload_8_sqIdx_flag | io_read_0_addr[9] &
    payload_9_sqIdx_flag | io_read_0_addr[10] & payload_10_sqIdx_flag | io_read_0_addr[11] & payload_11_sqIdx_flag |
    io_read_0_addr[12] & payload_12_sqIdx_flag | io_read_0_addr[13] & payload_13_sqIdx_flag | io_read_0_addr[14] &
    payload_14_sqIdx_flag | _io_read_0_data_T_403; // @[Mux.scala 27:73]
  assign io_read_0_data_sqIdx_value = _io_read_0_data_T_386 | _io_read_0_data_T_372; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_foldpc = _io_read_1_data_T_3300 | _io_read_1_data_T_3286; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_trigger_backendEn_0 = io_read_1_addr[0] & payload_0_cf_trigger_backendEn_0 | io_read_1_addr[1
    ] & payload_1_cf_trigger_backendEn_0 | io_read_1_addr[2] & payload_2_cf_trigger_backendEn_0 | io_read_1_addr[3] &
    payload_3_cf_trigger_backendEn_0 | io_read_1_addr[4] & payload_4_cf_trigger_backendEn_0 | io_read_1_addr[5] &
    payload_5_cf_trigger_backendEn_0 | io_read_1_addr[6] & payload_6_cf_trigger_backendEn_0 | io_read_1_addr[7] &
    payload_7_cf_trigger_backendEn_0 | io_read_1_addr[8] & payload_8_cf_trigger_backendEn_0 | io_read_1_addr[9] &
    payload_9_cf_trigger_backendEn_0 | io_read_1_addr[10] & payload_10_cf_trigger_backendEn_0 | io_read_1_addr[11] &
    payload_11_cf_trigger_backendEn_0 | io_read_1_addr[12] & payload_12_cf_trigger_backendEn_0 | io_read_1_addr[13] &
    payload_13_cf_trigger_backendEn_0 | io_read_1_addr[14] & payload_14_cf_trigger_backendEn_0 | _io_read_1_data_T_2604; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_trigger_backendEn_1 = io_read_1_addr[0] & payload_0_cf_trigger_backendEn_1 | io_read_1_addr[1
    ] & payload_1_cf_trigger_backendEn_1 | io_read_1_addr[2] & payload_2_cf_trigger_backendEn_1 | io_read_1_addr[3] &
    payload_3_cf_trigger_backendEn_1 | io_read_1_addr[4] & payload_4_cf_trigger_backendEn_1 | io_read_1_addr[5] &
    payload_5_cf_trigger_backendEn_1 | io_read_1_addr[6] & payload_6_cf_trigger_backendEn_1 | io_read_1_addr[7] &
    payload_7_cf_trigger_backendEn_1 | io_read_1_addr[8] & payload_8_cf_trigger_backendEn_1 | io_read_1_addr[9] &
    payload_9_cf_trigger_backendEn_1 | io_read_1_addr[10] & payload_10_cf_trigger_backendEn_1 | io_read_1_addr[11] &
    payload_11_cf_trigger_backendEn_1 | io_read_1_addr[12] & payload_12_cf_trigger_backendEn_1 | io_read_1_addr[13] &
    payload_13_cf_trigger_backendEn_1 | io_read_1_addr[14] & payload_14_cf_trigger_backendEn_1 | _io_read_1_data_T_2635; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pd_isRVC = io_read_1_addr[0] & payload_0_cf_pd_isRVC | io_read_1_addr[1] &
    payload_1_cf_pd_isRVC | io_read_1_addr[2] & payload_2_cf_pd_isRVC | io_read_1_addr[3] & payload_3_cf_pd_isRVC |
    io_read_1_addr[4] & payload_4_cf_pd_isRVC | io_read_1_addr[5] & payload_5_cf_pd_isRVC | io_read_1_addr[6] &
    payload_6_cf_pd_isRVC | io_read_1_addr[7] & payload_7_cf_pd_isRVC | io_read_1_addr[8] & payload_8_cf_pd_isRVC |
    io_read_1_addr[9] & payload_9_cf_pd_isRVC | io_read_1_addr[10] & payload_10_cf_pd_isRVC | io_read_1_addr[11] &
    payload_11_cf_pd_isRVC | io_read_1_addr[12] & payload_12_cf_pd_isRVC | io_read_1_addr[13] & payload_13_cf_pd_isRVC
     | io_read_1_addr[14] & payload_14_cf_pd_isRVC | _io_read_1_data_T_2356; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pd_brType = _io_read_1_data_T_2339 | _io_read_1_data_T_2325; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pd_isCall = io_read_1_addr[0] & payload_0_cf_pd_isCall | io_read_1_addr[1] &
    payload_1_cf_pd_isCall | io_read_1_addr[2] & payload_2_cf_pd_isCall | io_read_1_addr[3] & payload_3_cf_pd_isCall |
    io_read_1_addr[4] & payload_4_cf_pd_isCall | io_read_1_addr[5] & payload_5_cf_pd_isCall | io_read_1_addr[6] &
    payload_6_cf_pd_isCall | io_read_1_addr[7] & payload_7_cf_pd_isCall | io_read_1_addr[8] & payload_8_cf_pd_isCall |
    io_read_1_addr[9] & payload_9_cf_pd_isCall | io_read_1_addr[10] & payload_10_cf_pd_isCall | io_read_1_addr[11] &
    payload_11_cf_pd_isCall | io_read_1_addr[12] & payload_12_cf_pd_isCall | io_read_1_addr[13] &
    payload_13_cf_pd_isCall | io_read_1_addr[14] & payload_14_cf_pd_isCall | _io_read_1_data_T_2294; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pd_isRet = io_read_1_addr[0] & payload_0_cf_pd_isRet | io_read_1_addr[1] &
    payload_1_cf_pd_isRet | io_read_1_addr[2] & payload_2_cf_pd_isRet | io_read_1_addr[3] & payload_3_cf_pd_isRet |
    io_read_1_addr[4] & payload_4_cf_pd_isRet | io_read_1_addr[5] & payload_5_cf_pd_isRet | io_read_1_addr[6] &
    payload_6_cf_pd_isRet | io_read_1_addr[7] & payload_7_cf_pd_isRet | io_read_1_addr[8] & payload_8_cf_pd_isRet |
    io_read_1_addr[9] & payload_9_cf_pd_isRet | io_read_1_addr[10] & payload_10_cf_pd_isRet | io_read_1_addr[11] &
    payload_11_cf_pd_isRet | io_read_1_addr[12] & payload_12_cf_pd_isRet | io_read_1_addr[13] & payload_13_cf_pd_isRet
     | io_read_1_addr[14] & payload_14_cf_pd_isRet | _io_read_1_data_T_2263; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pred_taken = io_read_1_addr[0] & payload_0_cf_pred_taken | io_read_1_addr[1] &
    payload_1_cf_pred_taken | io_read_1_addr[2] & payload_2_cf_pred_taken | io_read_1_addr[3] & payload_3_cf_pred_taken
     | io_read_1_addr[4] & payload_4_cf_pred_taken | io_read_1_addr[5] & payload_5_cf_pred_taken | io_read_1_addr[6] &
    payload_6_cf_pred_taken | io_read_1_addr[7] & payload_7_cf_pred_taken | io_read_1_addr[8] & payload_8_cf_pred_taken
     | io_read_1_addr[9] & payload_9_cf_pred_taken | io_read_1_addr[10] & payload_10_cf_pred_taken | io_read_1_addr[11]
     & payload_11_cf_pred_taken | io_read_1_addr[12] & payload_12_cf_pred_taken | io_read_1_addr[13] &
    payload_13_cf_pred_taken | io_read_1_addr[14] & payload_14_cf_pred_taken | _io_read_1_data_T_2232; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_storeSetHit = io_read_1_addr[0] & payload_0_cf_storeSetHit | io_read_1_addr[1] &
    payload_1_cf_storeSetHit | io_read_1_addr[2] & payload_2_cf_storeSetHit | io_read_1_addr[3] &
    payload_3_cf_storeSetHit | io_read_1_addr[4] & payload_4_cf_storeSetHit | io_read_1_addr[5] &
    payload_5_cf_storeSetHit | io_read_1_addr[6] & payload_6_cf_storeSetHit | io_read_1_addr[7] &
    payload_7_cf_storeSetHit | io_read_1_addr[8] & payload_8_cf_storeSetHit | io_read_1_addr[9] &
    payload_9_cf_storeSetHit | io_read_1_addr[10] & payload_10_cf_storeSetHit | io_read_1_addr[11] &
    payload_11_cf_storeSetHit | io_read_1_addr[12] & payload_12_cf_storeSetHit | io_read_1_addr[13] &
    payload_13_cf_storeSetHit | io_read_1_addr[14] & payload_14_cf_storeSetHit | _io_read_1_data_T_2170; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_waitForRobIdx_flag = io_read_1_addr[0] & payload_0_cf_waitForRobIdx_flag | io_read_1_addr[1]
     & payload_1_cf_waitForRobIdx_flag | io_read_1_addr[2] & payload_2_cf_waitForRobIdx_flag | io_read_1_addr[3] &
    payload_3_cf_waitForRobIdx_flag | io_read_1_addr[4] & payload_4_cf_waitForRobIdx_flag | io_read_1_addr[5] &
    payload_5_cf_waitForRobIdx_flag | io_read_1_addr[6] & payload_6_cf_waitForRobIdx_flag | io_read_1_addr[7] &
    payload_7_cf_waitForRobIdx_flag | io_read_1_addr[8] & payload_8_cf_waitForRobIdx_flag | io_read_1_addr[9] &
    payload_9_cf_waitForRobIdx_flag | io_read_1_addr[10] & payload_10_cf_waitForRobIdx_flag | io_read_1_addr[11] &
    payload_11_cf_waitForRobIdx_flag | io_read_1_addr[12] & payload_12_cf_waitForRobIdx_flag | io_read_1_addr[13] &
    payload_13_cf_waitForRobIdx_flag | io_read_1_addr[14] & payload_14_cf_waitForRobIdx_flag | _io_read_1_data_T_2139; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_waitForRobIdx_value = _io_read_1_data_T_2122 | _io_read_1_data_T_2108; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_loadWaitBit = io_read_1_addr[0] & payload_0_cf_loadWaitBit | io_read_1_addr[1] &
    payload_1_cf_loadWaitBit | io_read_1_addr[2] & payload_2_cf_loadWaitBit | io_read_1_addr[3] &
    payload_3_cf_loadWaitBit | io_read_1_addr[4] & payload_4_cf_loadWaitBit | io_read_1_addr[5] &
    payload_5_cf_loadWaitBit | io_read_1_addr[6] & payload_6_cf_loadWaitBit | io_read_1_addr[7] &
    payload_7_cf_loadWaitBit | io_read_1_addr[8] & payload_8_cf_loadWaitBit | io_read_1_addr[9] &
    payload_9_cf_loadWaitBit | io_read_1_addr[10] & payload_10_cf_loadWaitBit | io_read_1_addr[11] &
    payload_11_cf_loadWaitBit | io_read_1_addr[12] & payload_12_cf_loadWaitBit | io_read_1_addr[13] &
    payload_13_cf_loadWaitBit | io_read_1_addr[14] & payload_14_cf_loadWaitBit | _io_read_1_data_T_2077; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_loadWaitStrict = io_read_1_addr[0] & payload_0_cf_loadWaitStrict | io_read_1_addr[1] &
    payload_1_cf_loadWaitStrict | io_read_1_addr[2] & payload_2_cf_loadWaitStrict | io_read_1_addr[3] &
    payload_3_cf_loadWaitStrict | io_read_1_addr[4] & payload_4_cf_loadWaitStrict | io_read_1_addr[5] &
    payload_5_cf_loadWaitStrict | io_read_1_addr[6] & payload_6_cf_loadWaitStrict | io_read_1_addr[7] &
    payload_7_cf_loadWaitStrict | io_read_1_addr[8] & payload_8_cf_loadWaitStrict | io_read_1_addr[9] &
    payload_9_cf_loadWaitStrict | io_read_1_addr[10] & payload_10_cf_loadWaitStrict | io_read_1_addr[11] &
    payload_11_cf_loadWaitStrict | io_read_1_addr[12] & payload_12_cf_loadWaitStrict | io_read_1_addr[13] &
    payload_13_cf_loadWaitStrict | io_read_1_addr[14] & payload_14_cf_loadWaitStrict | _io_read_1_data_T_2046; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_ssid = _io_read_1_data_T_2029 | _io_read_1_data_T_2015; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_ftqPtr_flag = io_read_1_addr[0] & payload_0_cf_ftqPtr_flag | io_read_1_addr[1] &
    payload_1_cf_ftqPtr_flag | io_read_1_addr[2] & payload_2_cf_ftqPtr_flag | io_read_1_addr[3] &
    payload_3_cf_ftqPtr_flag | io_read_1_addr[4] & payload_4_cf_ftqPtr_flag | io_read_1_addr[5] &
    payload_5_cf_ftqPtr_flag | io_read_1_addr[6] & payload_6_cf_ftqPtr_flag | io_read_1_addr[7] &
    payload_7_cf_ftqPtr_flag | io_read_1_addr[8] & payload_8_cf_ftqPtr_flag | io_read_1_addr[9] &
    payload_9_cf_ftqPtr_flag | io_read_1_addr[10] & payload_10_cf_ftqPtr_flag | io_read_1_addr[11] &
    payload_11_cf_ftqPtr_flag | io_read_1_addr[12] & payload_12_cf_ftqPtr_flag | io_read_1_addr[13] &
    payload_13_cf_ftqPtr_flag | io_read_1_addr[14] & payload_14_cf_ftqPtr_flag | _io_read_1_data_T_1984; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_ftqPtr_value = _io_read_1_data_T_1967 | _io_read_1_data_T_1953; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_ftqOffset = _io_read_1_data_T_1936 | _io_read_1_data_T_1922; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fuType = _io_read_1_data_T_1657 | _io_read_1_data_T_1643; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fuOpType = _io_read_1_data_T_1626 | _io_read_1_data_T_1612; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_rfWen = io_read_1_addr[0] & payload_0_ctrl_rfWen | io_read_1_addr[1] & payload_1_ctrl_rfWen
     | io_read_1_addr[2] & payload_2_ctrl_rfWen | io_read_1_addr[3] & payload_3_ctrl_rfWen | io_read_1_addr[4] &
    payload_4_ctrl_rfWen | io_read_1_addr[5] & payload_5_ctrl_rfWen | io_read_1_addr[6] & payload_6_ctrl_rfWen |
    io_read_1_addr[7] & payload_7_ctrl_rfWen | io_read_1_addr[8] & payload_8_ctrl_rfWen | io_read_1_addr[9] &
    payload_9_ctrl_rfWen | io_read_1_addr[10] & payload_10_ctrl_rfWen | io_read_1_addr[11] & payload_11_ctrl_rfWen |
    io_read_1_addr[12] & payload_12_ctrl_rfWen | io_read_1_addr[13] & payload_13_ctrl_rfWen | io_read_1_addr[14] &
    payload_14_ctrl_rfWen | _io_read_1_data_T_1581; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpWen = io_read_1_addr[0] & payload_0_ctrl_fpWen | io_read_1_addr[1] & payload_1_ctrl_fpWen
     | io_read_1_addr[2] & payload_2_ctrl_fpWen | io_read_1_addr[3] & payload_3_ctrl_fpWen | io_read_1_addr[4] &
    payload_4_ctrl_fpWen | io_read_1_addr[5] & payload_5_ctrl_fpWen | io_read_1_addr[6] & payload_6_ctrl_fpWen |
    io_read_1_addr[7] & payload_7_ctrl_fpWen | io_read_1_addr[8] & payload_8_ctrl_fpWen | io_read_1_addr[9] &
    payload_9_ctrl_fpWen | io_read_1_addr[10] & payload_10_ctrl_fpWen | io_read_1_addr[11] & payload_11_ctrl_fpWen |
    io_read_1_addr[12] & payload_12_ctrl_fpWen | io_read_1_addr[13] & payload_13_ctrl_fpWen | io_read_1_addr[14] &
    payload_14_ctrl_fpWen | _io_read_1_data_T_1550; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_imm = _io_read_1_data_T_1378 | _io_read_1_data_T_1364; // @[Mux.scala 27:73]
  assign io_read_1_data_pdest = _io_read_1_data_T_603 | _io_read_1_data_T_589; // @[Mux.scala 27:73]
  assign io_read_1_data_robIdx_flag = io_read_1_addr[0] & payload_0_robIdx_flag | io_read_1_addr[1] &
    payload_1_robIdx_flag | io_read_1_addr[2] & payload_2_robIdx_flag | io_read_1_addr[3] & payload_3_robIdx_flag |
    io_read_1_addr[4] & payload_4_robIdx_flag | io_read_1_addr[5] & payload_5_robIdx_flag | io_read_1_addr[6] &
    payload_6_robIdx_flag | io_read_1_addr[7] & payload_7_robIdx_flag | io_read_1_addr[8] & payload_8_robIdx_flag |
    io_read_1_addr[9] & payload_9_robIdx_flag | io_read_1_addr[10] & payload_10_robIdx_flag | io_read_1_addr[11] &
    payload_11_robIdx_flag | io_read_1_addr[12] & payload_12_robIdx_flag | io_read_1_addr[13] & payload_13_robIdx_flag
     | io_read_1_addr[14] & payload_14_robIdx_flag | _io_read_1_data_T_527; // @[Mux.scala 27:73]
  assign io_read_1_data_robIdx_value = _io_read_1_data_T_510 | _io_read_1_data_T_496; // @[Mux.scala 27:73]
  assign io_read_1_data_lqIdx_flag = io_read_1_addr[0] & payload_0_lqIdx_flag | io_read_1_addr[1] & payload_1_lqIdx_flag
     | io_read_1_addr[2] & payload_2_lqIdx_flag | io_read_1_addr[3] & payload_3_lqIdx_flag | io_read_1_addr[4] &
    payload_4_lqIdx_flag | io_read_1_addr[5] & payload_5_lqIdx_flag | io_read_1_addr[6] & payload_6_lqIdx_flag |
    io_read_1_addr[7] & payload_7_lqIdx_flag | io_read_1_addr[8] & payload_8_lqIdx_flag | io_read_1_addr[9] &
    payload_9_lqIdx_flag | io_read_1_addr[10] & payload_10_lqIdx_flag | io_read_1_addr[11] & payload_11_lqIdx_flag |
    io_read_1_addr[12] & payload_12_lqIdx_flag | io_read_1_addr[13] & payload_13_lqIdx_flag | io_read_1_addr[14] &
    payload_14_lqIdx_flag | _io_read_1_data_T_465; // @[Mux.scala 27:73]
  assign io_read_1_data_lqIdx_value = _io_read_1_data_T_448 | _io_read_1_data_T_434; // @[Mux.scala 27:73]
  assign io_read_1_data_sqIdx_flag = io_read_1_addr[0] & payload_0_sqIdx_flag | io_read_1_addr[1] & payload_1_sqIdx_flag
     | io_read_1_addr[2] & payload_2_sqIdx_flag | io_read_1_addr[3] & payload_3_sqIdx_flag | io_read_1_addr[4] &
    payload_4_sqIdx_flag | io_read_1_addr[5] & payload_5_sqIdx_flag | io_read_1_addr[6] & payload_6_sqIdx_flag |
    io_read_1_addr[7] & payload_7_sqIdx_flag | io_read_1_addr[8] & payload_8_sqIdx_flag | io_read_1_addr[9] &
    payload_9_sqIdx_flag | io_read_1_addr[10] & payload_10_sqIdx_flag | io_read_1_addr[11] & payload_11_sqIdx_flag |
    io_read_1_addr[12] & payload_12_sqIdx_flag | io_read_1_addr[13] & payload_13_sqIdx_flag | io_read_1_addr[14] &
    payload_14_sqIdx_flag | _io_read_1_data_T_403; // @[Mux.scala 27:73]
  assign io_read_1_data_sqIdx_value = _io_read_1_data_T_386 | _io_read_1_data_T_372; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_foldpc = _io_read_2_data_T_3300 | _io_read_2_data_T_3286; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_trigger_backendEn_0 = io_read_2_addr[0] & payload_0_cf_trigger_backendEn_0 | io_read_2_addr[1
    ] & payload_1_cf_trigger_backendEn_0 | io_read_2_addr[2] & payload_2_cf_trigger_backendEn_0 | io_read_2_addr[3] &
    payload_3_cf_trigger_backendEn_0 | io_read_2_addr[4] & payload_4_cf_trigger_backendEn_0 | io_read_2_addr[5] &
    payload_5_cf_trigger_backendEn_0 | io_read_2_addr[6] & payload_6_cf_trigger_backendEn_0 | io_read_2_addr[7] &
    payload_7_cf_trigger_backendEn_0 | io_read_2_addr[8] & payload_8_cf_trigger_backendEn_0 | io_read_2_addr[9] &
    payload_9_cf_trigger_backendEn_0 | io_read_2_addr[10] & payload_10_cf_trigger_backendEn_0 | io_read_2_addr[11] &
    payload_11_cf_trigger_backendEn_0 | io_read_2_addr[12] & payload_12_cf_trigger_backendEn_0 | io_read_2_addr[13] &
    payload_13_cf_trigger_backendEn_0 | io_read_2_addr[14] & payload_14_cf_trigger_backendEn_0 | _io_read_2_data_T_2604; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_trigger_backendEn_1 = io_read_2_addr[0] & payload_0_cf_trigger_backendEn_1 | io_read_2_addr[1
    ] & payload_1_cf_trigger_backendEn_1 | io_read_2_addr[2] & payload_2_cf_trigger_backendEn_1 | io_read_2_addr[3] &
    payload_3_cf_trigger_backendEn_1 | io_read_2_addr[4] & payload_4_cf_trigger_backendEn_1 | io_read_2_addr[5] &
    payload_5_cf_trigger_backendEn_1 | io_read_2_addr[6] & payload_6_cf_trigger_backendEn_1 | io_read_2_addr[7] &
    payload_7_cf_trigger_backendEn_1 | io_read_2_addr[8] & payload_8_cf_trigger_backendEn_1 | io_read_2_addr[9] &
    payload_9_cf_trigger_backendEn_1 | io_read_2_addr[10] & payload_10_cf_trigger_backendEn_1 | io_read_2_addr[11] &
    payload_11_cf_trigger_backendEn_1 | io_read_2_addr[12] & payload_12_cf_trigger_backendEn_1 | io_read_2_addr[13] &
    payload_13_cf_trigger_backendEn_1 | io_read_2_addr[14] & payload_14_cf_trigger_backendEn_1 | _io_read_2_data_T_2635; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_pd_isRVC = io_read_2_addr[0] & payload_0_cf_pd_isRVC | io_read_2_addr[1] &
    payload_1_cf_pd_isRVC | io_read_2_addr[2] & payload_2_cf_pd_isRVC | io_read_2_addr[3] & payload_3_cf_pd_isRVC |
    io_read_2_addr[4] & payload_4_cf_pd_isRVC | io_read_2_addr[5] & payload_5_cf_pd_isRVC | io_read_2_addr[6] &
    payload_6_cf_pd_isRVC | io_read_2_addr[7] & payload_7_cf_pd_isRVC | io_read_2_addr[8] & payload_8_cf_pd_isRVC |
    io_read_2_addr[9] & payload_9_cf_pd_isRVC | io_read_2_addr[10] & payload_10_cf_pd_isRVC | io_read_2_addr[11] &
    payload_11_cf_pd_isRVC | io_read_2_addr[12] & payload_12_cf_pd_isRVC | io_read_2_addr[13] & payload_13_cf_pd_isRVC
     | io_read_2_addr[14] & payload_14_cf_pd_isRVC | _io_read_2_data_T_2356; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_pd_brType = _io_read_2_data_T_2339 | _io_read_2_data_T_2325; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_pd_isCall = io_read_2_addr[0] & payload_0_cf_pd_isCall | io_read_2_addr[1] &
    payload_1_cf_pd_isCall | io_read_2_addr[2] & payload_2_cf_pd_isCall | io_read_2_addr[3] & payload_3_cf_pd_isCall |
    io_read_2_addr[4] & payload_4_cf_pd_isCall | io_read_2_addr[5] & payload_5_cf_pd_isCall | io_read_2_addr[6] &
    payload_6_cf_pd_isCall | io_read_2_addr[7] & payload_7_cf_pd_isCall | io_read_2_addr[8] & payload_8_cf_pd_isCall |
    io_read_2_addr[9] & payload_9_cf_pd_isCall | io_read_2_addr[10] & payload_10_cf_pd_isCall | io_read_2_addr[11] &
    payload_11_cf_pd_isCall | io_read_2_addr[12] & payload_12_cf_pd_isCall | io_read_2_addr[13] &
    payload_13_cf_pd_isCall | io_read_2_addr[14] & payload_14_cf_pd_isCall | _io_read_2_data_T_2294; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_pd_isRet = io_read_2_addr[0] & payload_0_cf_pd_isRet | io_read_2_addr[1] &
    payload_1_cf_pd_isRet | io_read_2_addr[2] & payload_2_cf_pd_isRet | io_read_2_addr[3] & payload_3_cf_pd_isRet |
    io_read_2_addr[4] & payload_4_cf_pd_isRet | io_read_2_addr[5] & payload_5_cf_pd_isRet | io_read_2_addr[6] &
    payload_6_cf_pd_isRet | io_read_2_addr[7] & payload_7_cf_pd_isRet | io_read_2_addr[8] & payload_8_cf_pd_isRet |
    io_read_2_addr[9] & payload_9_cf_pd_isRet | io_read_2_addr[10] & payload_10_cf_pd_isRet | io_read_2_addr[11] &
    payload_11_cf_pd_isRet | io_read_2_addr[12] & payload_12_cf_pd_isRet | io_read_2_addr[13] & payload_13_cf_pd_isRet
     | io_read_2_addr[14] & payload_14_cf_pd_isRet | _io_read_2_data_T_2263; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_pred_taken = io_read_2_addr[0] & payload_0_cf_pred_taken | io_read_2_addr[1] &
    payload_1_cf_pred_taken | io_read_2_addr[2] & payload_2_cf_pred_taken | io_read_2_addr[3] & payload_3_cf_pred_taken
     | io_read_2_addr[4] & payload_4_cf_pred_taken | io_read_2_addr[5] & payload_5_cf_pred_taken | io_read_2_addr[6] &
    payload_6_cf_pred_taken | io_read_2_addr[7] & payload_7_cf_pred_taken | io_read_2_addr[8] & payload_8_cf_pred_taken
     | io_read_2_addr[9] & payload_9_cf_pred_taken | io_read_2_addr[10] & payload_10_cf_pred_taken | io_read_2_addr[11]
     & payload_11_cf_pred_taken | io_read_2_addr[12] & payload_12_cf_pred_taken | io_read_2_addr[13] &
    payload_13_cf_pred_taken | io_read_2_addr[14] & payload_14_cf_pred_taken | _io_read_2_data_T_2232; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_storeSetHit = io_read_2_addr[0] & payload_0_cf_storeSetHit | io_read_2_addr[1] &
    payload_1_cf_storeSetHit | io_read_2_addr[2] & payload_2_cf_storeSetHit | io_read_2_addr[3] &
    payload_3_cf_storeSetHit | io_read_2_addr[4] & payload_4_cf_storeSetHit | io_read_2_addr[5] &
    payload_5_cf_storeSetHit | io_read_2_addr[6] & payload_6_cf_storeSetHit | io_read_2_addr[7] &
    payload_7_cf_storeSetHit | io_read_2_addr[8] & payload_8_cf_storeSetHit | io_read_2_addr[9] &
    payload_9_cf_storeSetHit | io_read_2_addr[10] & payload_10_cf_storeSetHit | io_read_2_addr[11] &
    payload_11_cf_storeSetHit | io_read_2_addr[12] & payload_12_cf_storeSetHit | io_read_2_addr[13] &
    payload_13_cf_storeSetHit | io_read_2_addr[14] & payload_14_cf_storeSetHit | _io_read_2_data_T_2170; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_waitForRobIdx_flag = io_read_2_addr[0] & payload_0_cf_waitForRobIdx_flag | io_read_2_addr[1]
     & payload_1_cf_waitForRobIdx_flag | io_read_2_addr[2] & payload_2_cf_waitForRobIdx_flag | io_read_2_addr[3] &
    payload_3_cf_waitForRobIdx_flag | io_read_2_addr[4] & payload_4_cf_waitForRobIdx_flag | io_read_2_addr[5] &
    payload_5_cf_waitForRobIdx_flag | io_read_2_addr[6] & payload_6_cf_waitForRobIdx_flag | io_read_2_addr[7] &
    payload_7_cf_waitForRobIdx_flag | io_read_2_addr[8] & payload_8_cf_waitForRobIdx_flag | io_read_2_addr[9] &
    payload_9_cf_waitForRobIdx_flag | io_read_2_addr[10] & payload_10_cf_waitForRobIdx_flag | io_read_2_addr[11] &
    payload_11_cf_waitForRobIdx_flag | io_read_2_addr[12] & payload_12_cf_waitForRobIdx_flag | io_read_2_addr[13] &
    payload_13_cf_waitForRobIdx_flag | io_read_2_addr[14] & payload_14_cf_waitForRobIdx_flag | _io_read_2_data_T_2139; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_waitForRobIdx_value = _io_read_2_data_T_2122 | _io_read_2_data_T_2108; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_loadWaitBit = io_read_2_addr[0] & payload_0_cf_loadWaitBit | io_read_2_addr[1] &
    payload_1_cf_loadWaitBit | io_read_2_addr[2] & payload_2_cf_loadWaitBit | io_read_2_addr[3] &
    payload_3_cf_loadWaitBit | io_read_2_addr[4] & payload_4_cf_loadWaitBit | io_read_2_addr[5] &
    payload_5_cf_loadWaitBit | io_read_2_addr[6] & payload_6_cf_loadWaitBit | io_read_2_addr[7] &
    payload_7_cf_loadWaitBit | io_read_2_addr[8] & payload_8_cf_loadWaitBit | io_read_2_addr[9] &
    payload_9_cf_loadWaitBit | io_read_2_addr[10] & payload_10_cf_loadWaitBit | io_read_2_addr[11] &
    payload_11_cf_loadWaitBit | io_read_2_addr[12] & payload_12_cf_loadWaitBit | io_read_2_addr[13] &
    payload_13_cf_loadWaitBit | io_read_2_addr[14] & payload_14_cf_loadWaitBit | _io_read_2_data_T_2077; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_loadWaitStrict = io_read_2_addr[0] & payload_0_cf_loadWaitStrict | io_read_2_addr[1] &
    payload_1_cf_loadWaitStrict | io_read_2_addr[2] & payload_2_cf_loadWaitStrict | io_read_2_addr[3] &
    payload_3_cf_loadWaitStrict | io_read_2_addr[4] & payload_4_cf_loadWaitStrict | io_read_2_addr[5] &
    payload_5_cf_loadWaitStrict | io_read_2_addr[6] & payload_6_cf_loadWaitStrict | io_read_2_addr[7] &
    payload_7_cf_loadWaitStrict | io_read_2_addr[8] & payload_8_cf_loadWaitStrict | io_read_2_addr[9] &
    payload_9_cf_loadWaitStrict | io_read_2_addr[10] & payload_10_cf_loadWaitStrict | io_read_2_addr[11] &
    payload_11_cf_loadWaitStrict | io_read_2_addr[12] & payload_12_cf_loadWaitStrict | io_read_2_addr[13] &
    payload_13_cf_loadWaitStrict | io_read_2_addr[14] & payload_14_cf_loadWaitStrict | _io_read_2_data_T_2046; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_ssid = _io_read_2_data_T_2029 | _io_read_2_data_T_2015; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_ftqPtr_flag = io_read_2_addr[0] & payload_0_cf_ftqPtr_flag | io_read_2_addr[1] &
    payload_1_cf_ftqPtr_flag | io_read_2_addr[2] & payload_2_cf_ftqPtr_flag | io_read_2_addr[3] &
    payload_3_cf_ftqPtr_flag | io_read_2_addr[4] & payload_4_cf_ftqPtr_flag | io_read_2_addr[5] &
    payload_5_cf_ftqPtr_flag | io_read_2_addr[6] & payload_6_cf_ftqPtr_flag | io_read_2_addr[7] &
    payload_7_cf_ftqPtr_flag | io_read_2_addr[8] & payload_8_cf_ftqPtr_flag | io_read_2_addr[9] &
    payload_9_cf_ftqPtr_flag | io_read_2_addr[10] & payload_10_cf_ftqPtr_flag | io_read_2_addr[11] &
    payload_11_cf_ftqPtr_flag | io_read_2_addr[12] & payload_12_cf_ftqPtr_flag | io_read_2_addr[13] &
    payload_13_cf_ftqPtr_flag | io_read_2_addr[14] & payload_14_cf_ftqPtr_flag | _io_read_2_data_T_1984; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_ftqPtr_value = _io_read_2_data_T_1967 | _io_read_2_data_T_1953; // @[Mux.scala 27:73]
  assign io_read_2_data_cf_ftqOffset = _io_read_2_data_T_1936 | _io_read_2_data_T_1922; // @[Mux.scala 27:73]
  assign io_read_2_data_ctrl_fuType = _io_read_2_data_T_1657 | _io_read_2_data_T_1643; // @[Mux.scala 27:73]
  assign io_read_2_data_ctrl_fuOpType = _io_read_2_data_T_1626 | _io_read_2_data_T_1612; // @[Mux.scala 27:73]
  assign io_read_2_data_ctrl_rfWen = io_read_2_addr[0] & payload_0_ctrl_rfWen | io_read_2_addr[1] & payload_1_ctrl_rfWen
     | io_read_2_addr[2] & payload_2_ctrl_rfWen | io_read_2_addr[3] & payload_3_ctrl_rfWen | io_read_2_addr[4] &
    payload_4_ctrl_rfWen | io_read_2_addr[5] & payload_5_ctrl_rfWen | io_read_2_addr[6] & payload_6_ctrl_rfWen |
    io_read_2_addr[7] & payload_7_ctrl_rfWen | io_read_2_addr[8] & payload_8_ctrl_rfWen | io_read_2_addr[9] &
    payload_9_ctrl_rfWen | io_read_2_addr[10] & payload_10_ctrl_rfWen | io_read_2_addr[11] & payload_11_ctrl_rfWen |
    io_read_2_addr[12] & payload_12_ctrl_rfWen | io_read_2_addr[13] & payload_13_ctrl_rfWen | io_read_2_addr[14] &
    payload_14_ctrl_rfWen | _io_read_2_data_T_1581; // @[Mux.scala 27:73]
  assign io_read_2_data_ctrl_fpWen = io_read_2_addr[0] & payload_0_ctrl_fpWen | io_read_2_addr[1] & payload_1_ctrl_fpWen
     | io_read_2_addr[2] & payload_2_ctrl_fpWen | io_read_2_addr[3] & payload_3_ctrl_fpWen | io_read_2_addr[4] &
    payload_4_ctrl_fpWen | io_read_2_addr[5] & payload_5_ctrl_fpWen | io_read_2_addr[6] & payload_6_ctrl_fpWen |
    io_read_2_addr[7] & payload_7_ctrl_fpWen | io_read_2_addr[8] & payload_8_ctrl_fpWen | io_read_2_addr[9] &
    payload_9_ctrl_fpWen | io_read_2_addr[10] & payload_10_ctrl_fpWen | io_read_2_addr[11] & payload_11_ctrl_fpWen |
    io_read_2_addr[12] & payload_12_ctrl_fpWen | io_read_2_addr[13] & payload_13_ctrl_fpWen | io_read_2_addr[14] &
    payload_14_ctrl_fpWen | _io_read_2_data_T_1550; // @[Mux.scala 27:73]
  assign io_read_2_data_ctrl_imm = _io_read_2_data_T_1378 | _io_read_2_data_T_1364; // @[Mux.scala 27:73]
  assign io_read_2_data_pdest = _io_read_2_data_T_603 | _io_read_2_data_T_589; // @[Mux.scala 27:73]
  assign io_read_2_data_robIdx_flag = io_read_2_addr[0] & payload_0_robIdx_flag | io_read_2_addr[1] &
    payload_1_robIdx_flag | io_read_2_addr[2] & payload_2_robIdx_flag | io_read_2_addr[3] & payload_3_robIdx_flag |
    io_read_2_addr[4] & payload_4_robIdx_flag | io_read_2_addr[5] & payload_5_robIdx_flag | io_read_2_addr[6] &
    payload_6_robIdx_flag | io_read_2_addr[7] & payload_7_robIdx_flag | io_read_2_addr[8] & payload_8_robIdx_flag |
    io_read_2_addr[9] & payload_9_robIdx_flag | io_read_2_addr[10] & payload_10_robIdx_flag | io_read_2_addr[11] &
    payload_11_robIdx_flag | io_read_2_addr[12] & payload_12_robIdx_flag | io_read_2_addr[13] & payload_13_robIdx_flag
     | io_read_2_addr[14] & payload_14_robIdx_flag | _io_read_2_data_T_527; // @[Mux.scala 27:73]
  assign io_read_2_data_robIdx_value = _io_read_2_data_T_510 | _io_read_2_data_T_496; // @[Mux.scala 27:73]
  assign io_read_2_data_lqIdx_flag = io_read_2_addr[0] & payload_0_lqIdx_flag | io_read_2_addr[1] & payload_1_lqIdx_flag
     | io_read_2_addr[2] & payload_2_lqIdx_flag | io_read_2_addr[3] & payload_3_lqIdx_flag | io_read_2_addr[4] &
    payload_4_lqIdx_flag | io_read_2_addr[5] & payload_5_lqIdx_flag | io_read_2_addr[6] & payload_6_lqIdx_flag |
    io_read_2_addr[7] & payload_7_lqIdx_flag | io_read_2_addr[8] & payload_8_lqIdx_flag | io_read_2_addr[9] &
    payload_9_lqIdx_flag | io_read_2_addr[10] & payload_10_lqIdx_flag | io_read_2_addr[11] & payload_11_lqIdx_flag |
    io_read_2_addr[12] & payload_12_lqIdx_flag | io_read_2_addr[13] & payload_13_lqIdx_flag | io_read_2_addr[14] &
    payload_14_lqIdx_flag | _io_read_2_data_T_465; // @[Mux.scala 27:73]
  assign io_read_2_data_lqIdx_value = _io_read_2_data_T_448 | _io_read_2_data_T_434; // @[Mux.scala 27:73]
  assign io_read_2_data_sqIdx_flag = io_read_2_addr[0] & payload_0_sqIdx_flag | io_read_2_addr[1] & payload_1_sqIdx_flag
     | io_read_2_addr[2] & payload_2_sqIdx_flag | io_read_2_addr[3] & payload_3_sqIdx_flag | io_read_2_addr[4] &
    payload_4_sqIdx_flag | io_read_2_addr[5] & payload_5_sqIdx_flag | io_read_2_addr[6] & payload_6_sqIdx_flag |
    io_read_2_addr[7] & payload_7_sqIdx_flag | io_read_2_addr[8] & payload_8_sqIdx_flag | io_read_2_addr[9] &
    payload_9_sqIdx_flag | io_read_2_addr[10] & payload_10_sqIdx_flag | io_read_2_addr[11] & payload_11_sqIdx_flag |
    io_read_2_addr[12] & payload_12_sqIdx_flag | io_read_2_addr[13] & payload_13_sqIdx_flag | io_read_2_addr[14] &
    payload_14_sqIdx_flag | _io_read_2_data_T_403; // @[Mux.scala 27:73]
  assign io_read_2_data_sqIdx_value = _io_read_2_data_T_386 | _io_read_2_data_T_372; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_foldpc <= wdata_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_trigger_backendEn_0 <= wdata_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_trigger_backendEn_1 <= wdata_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pd_isRVC <= wdata_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pd_brType <= wdata_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pd_isCall <= wdata_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pd_isRet <= wdata_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pred_taken <= wdata_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_storeSetHit <= wdata_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_waitForRobIdx_flag <= wdata_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_waitForRobIdx_value <= wdata_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_loadWaitBit <= wdata_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_loadWaitStrict <= wdata_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_ssid <= wdata_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_ftqPtr_flag <= wdata_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_ftqPtr_value <= wdata_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_ftqOffset <= wdata_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fuType <= wdata_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fuOpType <= wdata_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_rfWen <= wdata_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpWen <= wdata_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_imm <= wdata_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_pdest <= wdata_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_robIdx_flag <= wdata_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_robIdx_value <= wdata_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_lqIdx_flag <= wdata_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_lqIdx_value <= wdata_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_sqIdx_flag <= wdata_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_sqIdx_value <= wdata_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_foldpc <= wdata_1_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_trigger_backendEn_0 <= wdata_1_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_trigger_backendEn_1 <= wdata_1_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pd_isRVC <= wdata_1_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pd_brType <= wdata_1_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pd_isCall <= wdata_1_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pd_isRet <= wdata_1_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pred_taken <= wdata_1_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_storeSetHit <= wdata_1_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_waitForRobIdx_flag <= wdata_1_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_waitForRobIdx_value <= wdata_1_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_loadWaitBit <= wdata_1_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_loadWaitStrict <= wdata_1_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_ssid <= wdata_1_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_ftqPtr_flag <= wdata_1_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_ftqPtr_value <= wdata_1_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_ftqOffset <= wdata_1_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fuType <= wdata_1_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fuOpType <= wdata_1_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_rfWen <= wdata_1_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpWen <= wdata_1_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_imm <= wdata_1_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_pdest <= wdata_1_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_robIdx_flag <= wdata_1_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_robIdx_value <= wdata_1_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_lqIdx_flag <= wdata_1_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_lqIdx_value <= wdata_1_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_sqIdx_flag <= wdata_1_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_sqIdx_value <= wdata_1_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_foldpc <= wdata_2_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_trigger_backendEn_0 <= wdata_2_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_trigger_backendEn_1 <= wdata_2_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pd_isRVC <= wdata_2_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pd_brType <= wdata_2_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pd_isCall <= wdata_2_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pd_isRet <= wdata_2_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pred_taken <= wdata_2_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_storeSetHit <= wdata_2_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_waitForRobIdx_flag <= wdata_2_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_waitForRobIdx_value <= wdata_2_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_loadWaitBit <= wdata_2_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_loadWaitStrict <= wdata_2_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_ssid <= wdata_2_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_ftqPtr_flag <= wdata_2_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_ftqPtr_value <= wdata_2_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_ftqOffset <= wdata_2_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fuType <= wdata_2_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fuOpType <= wdata_2_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_rfWen <= wdata_2_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpWen <= wdata_2_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_imm <= wdata_2_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_pdest <= wdata_2_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_robIdx_flag <= wdata_2_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_robIdx_value <= wdata_2_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_lqIdx_flag <= wdata_2_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_lqIdx_value <= wdata_2_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_sqIdx_flag <= wdata_2_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_sqIdx_value <= wdata_2_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_foldpc <= wdata_3_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_trigger_backendEn_0 <= wdata_3_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_trigger_backendEn_1 <= wdata_3_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pd_isRVC <= wdata_3_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pd_brType <= wdata_3_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pd_isCall <= wdata_3_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pd_isRet <= wdata_3_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pred_taken <= wdata_3_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_storeSetHit <= wdata_3_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_waitForRobIdx_flag <= wdata_3_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_waitForRobIdx_value <= wdata_3_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_loadWaitBit <= wdata_3_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_loadWaitStrict <= wdata_3_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_ssid <= wdata_3_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_ftqPtr_flag <= wdata_3_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_ftqPtr_value <= wdata_3_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_ftqOffset <= wdata_3_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fuType <= wdata_3_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fuOpType <= wdata_3_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_rfWen <= wdata_3_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpWen <= wdata_3_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_imm <= wdata_3_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_pdest <= wdata_3_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_robIdx_flag <= wdata_3_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_robIdx_value <= wdata_3_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_lqIdx_flag <= wdata_3_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_lqIdx_value <= wdata_3_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_sqIdx_flag <= wdata_3_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_sqIdx_value <= wdata_3_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_foldpc <= wdata_4_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_trigger_backendEn_0 <= wdata_4_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_trigger_backendEn_1 <= wdata_4_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pd_isRVC <= wdata_4_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pd_brType <= wdata_4_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pd_isCall <= wdata_4_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pd_isRet <= wdata_4_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pred_taken <= wdata_4_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_storeSetHit <= wdata_4_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_waitForRobIdx_flag <= wdata_4_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_waitForRobIdx_value <= wdata_4_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_loadWaitBit <= wdata_4_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_loadWaitStrict <= wdata_4_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_ssid <= wdata_4_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_ftqPtr_flag <= wdata_4_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_ftqPtr_value <= wdata_4_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_ftqOffset <= wdata_4_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fuType <= wdata_4_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fuOpType <= wdata_4_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_rfWen <= wdata_4_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpWen <= wdata_4_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_imm <= wdata_4_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_pdest <= wdata_4_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_robIdx_flag <= wdata_4_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_robIdx_value <= wdata_4_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_lqIdx_flag <= wdata_4_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_lqIdx_value <= wdata_4_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_sqIdx_flag <= wdata_4_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_sqIdx_value <= wdata_4_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_foldpc <= wdata_5_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_trigger_backendEn_0 <= wdata_5_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_trigger_backendEn_1 <= wdata_5_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pd_isRVC <= wdata_5_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pd_brType <= wdata_5_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pd_isCall <= wdata_5_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pd_isRet <= wdata_5_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pred_taken <= wdata_5_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_storeSetHit <= wdata_5_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_waitForRobIdx_flag <= wdata_5_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_waitForRobIdx_value <= wdata_5_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_loadWaitBit <= wdata_5_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_loadWaitStrict <= wdata_5_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_ssid <= wdata_5_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_ftqPtr_flag <= wdata_5_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_ftqPtr_value <= wdata_5_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_ftqOffset <= wdata_5_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fuType <= wdata_5_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fuOpType <= wdata_5_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_rfWen <= wdata_5_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpWen <= wdata_5_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_imm <= wdata_5_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_pdest <= wdata_5_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_robIdx_flag <= wdata_5_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_robIdx_value <= wdata_5_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_lqIdx_flag <= wdata_5_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_lqIdx_value <= wdata_5_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_sqIdx_flag <= wdata_5_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_sqIdx_value <= wdata_5_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_foldpc <= wdata_6_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_trigger_backendEn_0 <= wdata_6_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_trigger_backendEn_1 <= wdata_6_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pd_isRVC <= wdata_6_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pd_brType <= wdata_6_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pd_isCall <= wdata_6_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pd_isRet <= wdata_6_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pred_taken <= wdata_6_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_storeSetHit <= wdata_6_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_waitForRobIdx_flag <= wdata_6_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_waitForRobIdx_value <= wdata_6_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_loadWaitBit <= wdata_6_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_loadWaitStrict <= wdata_6_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_ssid <= wdata_6_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_ftqPtr_flag <= wdata_6_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_ftqPtr_value <= wdata_6_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_ftqOffset <= wdata_6_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fuType <= wdata_6_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fuOpType <= wdata_6_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_rfWen <= wdata_6_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpWen <= wdata_6_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_imm <= wdata_6_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_pdest <= wdata_6_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_robIdx_flag <= wdata_6_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_robIdx_value <= wdata_6_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_lqIdx_flag <= wdata_6_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_lqIdx_value <= wdata_6_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_sqIdx_flag <= wdata_6_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_sqIdx_value <= wdata_6_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_foldpc <= wdata_7_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_trigger_backendEn_0 <= wdata_7_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_trigger_backendEn_1 <= wdata_7_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pd_isRVC <= wdata_7_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pd_brType <= wdata_7_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pd_isCall <= wdata_7_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pd_isRet <= wdata_7_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pred_taken <= wdata_7_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_storeSetHit <= wdata_7_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_waitForRobIdx_flag <= wdata_7_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_waitForRobIdx_value <= wdata_7_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_loadWaitBit <= wdata_7_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_loadWaitStrict <= wdata_7_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_ssid <= wdata_7_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_ftqPtr_flag <= wdata_7_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_ftqPtr_value <= wdata_7_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_ftqOffset <= wdata_7_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fuType <= wdata_7_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fuOpType <= wdata_7_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_rfWen <= wdata_7_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpWen <= wdata_7_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_imm <= wdata_7_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_pdest <= wdata_7_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_robIdx_flag <= wdata_7_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_robIdx_value <= wdata_7_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_lqIdx_flag <= wdata_7_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_lqIdx_value <= wdata_7_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_sqIdx_flag <= wdata_7_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_sqIdx_value <= wdata_7_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_foldpc <= wdata_8_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_trigger_backendEn_0 <= wdata_8_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_trigger_backendEn_1 <= wdata_8_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_pd_isRVC <= wdata_8_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_pd_brType <= wdata_8_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_pd_isCall <= wdata_8_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_pd_isRet <= wdata_8_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_pred_taken <= wdata_8_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_storeSetHit <= wdata_8_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_waitForRobIdx_flag <= wdata_8_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_waitForRobIdx_value <= wdata_8_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_loadWaitBit <= wdata_8_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_loadWaitStrict <= wdata_8_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_ssid <= wdata_8_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_ftqPtr_flag <= wdata_8_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_ftqPtr_value <= wdata_8_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_cf_ftqOffset <= wdata_8_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_ctrl_fuType <= wdata_8_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_ctrl_fuOpType <= wdata_8_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_ctrl_rfWen <= wdata_8_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_ctrl_fpWen <= wdata_8_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_ctrl_imm <= wdata_8_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_pdest <= wdata_8_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_robIdx_flag <= wdata_8_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_robIdx_value <= wdata_8_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_lqIdx_flag <= wdata_8_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_lqIdx_value <= wdata_8_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_sqIdx_flag <= wdata_8_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_8) begin // @[PayloadArray.scala 58:16]
      payload_8_sqIdx_value <= wdata_8_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_foldpc <= wdata_9_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_trigger_backendEn_0 <= wdata_9_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_trigger_backendEn_1 <= wdata_9_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_pd_isRVC <= wdata_9_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_pd_brType <= wdata_9_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_pd_isCall <= wdata_9_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_pd_isRet <= wdata_9_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_pred_taken <= wdata_9_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_storeSetHit <= wdata_9_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_waitForRobIdx_flag <= wdata_9_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_waitForRobIdx_value <= wdata_9_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_loadWaitBit <= wdata_9_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_loadWaitStrict <= wdata_9_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_ssid <= wdata_9_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_ftqPtr_flag <= wdata_9_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_ftqPtr_value <= wdata_9_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_cf_ftqOffset <= wdata_9_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_ctrl_fuType <= wdata_9_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_ctrl_fuOpType <= wdata_9_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_ctrl_rfWen <= wdata_9_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_ctrl_fpWen <= wdata_9_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_ctrl_imm <= wdata_9_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_pdest <= wdata_9_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_robIdx_flag <= wdata_9_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_robIdx_value <= wdata_9_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_lqIdx_flag <= wdata_9_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_lqIdx_value <= wdata_9_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_sqIdx_flag <= wdata_9_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_9) begin // @[PayloadArray.scala 58:16]
      payload_9_sqIdx_value <= wdata_9_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_foldpc <= wdata_10_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_trigger_backendEn_0 <= wdata_10_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_trigger_backendEn_1 <= wdata_10_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_pd_isRVC <= wdata_10_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_pd_brType <= wdata_10_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_pd_isCall <= wdata_10_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_pd_isRet <= wdata_10_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_pred_taken <= wdata_10_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_storeSetHit <= wdata_10_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_waitForRobIdx_flag <= wdata_10_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_waitForRobIdx_value <= wdata_10_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_loadWaitBit <= wdata_10_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_loadWaitStrict <= wdata_10_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_ssid <= wdata_10_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_ftqPtr_flag <= wdata_10_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_ftqPtr_value <= wdata_10_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_cf_ftqOffset <= wdata_10_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_ctrl_fuType <= wdata_10_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_ctrl_fuOpType <= wdata_10_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_ctrl_rfWen <= wdata_10_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_ctrl_fpWen <= wdata_10_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_ctrl_imm <= wdata_10_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_pdest <= wdata_10_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_robIdx_flag <= wdata_10_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_robIdx_value <= wdata_10_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_lqIdx_flag <= wdata_10_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_lqIdx_value <= wdata_10_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_sqIdx_flag <= wdata_10_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_10) begin // @[PayloadArray.scala 58:16]
      payload_10_sqIdx_value <= wdata_10_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_foldpc <= wdata_11_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_trigger_backendEn_0 <= wdata_11_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_trigger_backendEn_1 <= wdata_11_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_pd_isRVC <= wdata_11_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_pd_brType <= wdata_11_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_pd_isCall <= wdata_11_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_pd_isRet <= wdata_11_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_pred_taken <= wdata_11_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_storeSetHit <= wdata_11_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_waitForRobIdx_flag <= wdata_11_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_waitForRobIdx_value <= wdata_11_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_loadWaitBit <= wdata_11_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_loadWaitStrict <= wdata_11_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_ssid <= wdata_11_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_ftqPtr_flag <= wdata_11_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_ftqPtr_value <= wdata_11_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_cf_ftqOffset <= wdata_11_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_ctrl_fuType <= wdata_11_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_ctrl_fuOpType <= wdata_11_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_ctrl_rfWen <= wdata_11_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_ctrl_fpWen <= wdata_11_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_ctrl_imm <= wdata_11_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_pdest <= wdata_11_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_robIdx_flag <= wdata_11_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_robIdx_value <= wdata_11_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_lqIdx_flag <= wdata_11_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_lqIdx_value <= wdata_11_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_sqIdx_flag <= wdata_11_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_11) begin // @[PayloadArray.scala 58:16]
      payload_11_sqIdx_value <= wdata_11_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_foldpc <= wdata_12_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_trigger_backendEn_0 <= wdata_12_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_trigger_backendEn_1 <= wdata_12_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_pd_isRVC <= wdata_12_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_pd_brType <= wdata_12_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_pd_isCall <= wdata_12_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_pd_isRet <= wdata_12_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_pred_taken <= wdata_12_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_storeSetHit <= wdata_12_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_waitForRobIdx_flag <= wdata_12_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_waitForRobIdx_value <= wdata_12_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_loadWaitBit <= wdata_12_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_loadWaitStrict <= wdata_12_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_ssid <= wdata_12_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_ftqPtr_flag <= wdata_12_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_ftqPtr_value <= wdata_12_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_cf_ftqOffset <= wdata_12_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_ctrl_fuType <= wdata_12_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_ctrl_fuOpType <= wdata_12_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_ctrl_rfWen <= wdata_12_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_ctrl_fpWen <= wdata_12_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_ctrl_imm <= wdata_12_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_pdest <= wdata_12_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_robIdx_flag <= wdata_12_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_robIdx_value <= wdata_12_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_lqIdx_flag <= wdata_12_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_lqIdx_value <= wdata_12_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_sqIdx_flag <= wdata_12_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_12) begin // @[PayloadArray.scala 58:16]
      payload_12_sqIdx_value <= wdata_12_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_foldpc <= wdata_13_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_trigger_backendEn_0 <= wdata_13_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_trigger_backendEn_1 <= wdata_13_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_pd_isRVC <= wdata_13_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_pd_brType <= wdata_13_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_pd_isCall <= wdata_13_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_pd_isRet <= wdata_13_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_pred_taken <= wdata_13_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_storeSetHit <= wdata_13_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_waitForRobIdx_flag <= wdata_13_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_waitForRobIdx_value <= wdata_13_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_loadWaitBit <= wdata_13_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_loadWaitStrict <= wdata_13_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_ssid <= wdata_13_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_ftqPtr_flag <= wdata_13_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_ftqPtr_value <= wdata_13_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_cf_ftqOffset <= wdata_13_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_ctrl_fuType <= wdata_13_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_ctrl_fuOpType <= wdata_13_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_ctrl_rfWen <= wdata_13_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_ctrl_fpWen <= wdata_13_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_ctrl_imm <= wdata_13_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_pdest <= wdata_13_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_robIdx_flag <= wdata_13_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_robIdx_value <= wdata_13_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_lqIdx_flag <= wdata_13_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_lqIdx_value <= wdata_13_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_sqIdx_flag <= wdata_13_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_13) begin // @[PayloadArray.scala 58:16]
      payload_13_sqIdx_value <= wdata_13_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_foldpc <= wdata_14_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_trigger_backendEn_0 <= wdata_14_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_trigger_backendEn_1 <= wdata_14_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_pd_isRVC <= wdata_14_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_pd_brType <= wdata_14_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_pd_isCall <= wdata_14_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_pd_isRet <= wdata_14_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_pred_taken <= wdata_14_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_storeSetHit <= wdata_14_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_waitForRobIdx_flag <= wdata_14_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_waitForRobIdx_value <= wdata_14_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_loadWaitBit <= wdata_14_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_loadWaitStrict <= wdata_14_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_ssid <= wdata_14_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_ftqPtr_flag <= wdata_14_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_ftqPtr_value <= wdata_14_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_cf_ftqOffset <= wdata_14_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_ctrl_fuType <= wdata_14_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_ctrl_fuOpType <= wdata_14_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_ctrl_rfWen <= wdata_14_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_ctrl_fpWen <= wdata_14_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_ctrl_imm <= wdata_14_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_pdest <= wdata_14_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_robIdx_flag <= wdata_14_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_robIdx_value <= wdata_14_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_lqIdx_flag <= wdata_14_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_lqIdx_value <= wdata_14_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_sqIdx_flag <= wdata_14_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_14) begin // @[PayloadArray.scala 58:16]
      payload_14_sqIdx_value <= wdata_14_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_foldpc <= wdata_15_cf_foldpc; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_trigger_backendEn_0 <= wdata_15_cf_trigger_backendEn_0; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_trigger_backendEn_1 <= wdata_15_cf_trigger_backendEn_1; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_pd_isRVC <= wdata_15_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_pd_brType <= wdata_15_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_pd_isCall <= wdata_15_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_pd_isRet <= wdata_15_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_pred_taken <= wdata_15_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_storeSetHit <= wdata_15_cf_storeSetHit; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_waitForRobIdx_flag <= wdata_15_cf_waitForRobIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_waitForRobIdx_value <= wdata_15_cf_waitForRobIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_loadWaitBit <= wdata_15_cf_loadWaitBit; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_loadWaitStrict <= wdata_15_cf_loadWaitStrict; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_ssid <= wdata_15_cf_ssid; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_ftqPtr_flag <= wdata_15_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_ftqPtr_value <= wdata_15_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_cf_ftqOffset <= wdata_15_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_ctrl_fuType <= wdata_15_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_ctrl_fuOpType <= wdata_15_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_ctrl_rfWen <= wdata_15_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_ctrl_fpWen <= wdata_15_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_ctrl_imm <= wdata_15_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_pdest <= wdata_15_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_robIdx_flag <= wdata_15_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_robIdx_value <= wdata_15_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_lqIdx_flag <= wdata_15_lqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_lqIdx_value <= wdata_15_lqIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_sqIdx_flag <= wdata_15_sqIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_15) begin // @[PayloadArray.scala 58:16]
      payload_15_sqIdx_value <= wdata_15_sqIdx_value; // @[PayloadArray.scala 59:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  payload_0_cf_foldpc = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  payload_0_cf_trigger_backendEn_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  payload_0_cf_trigger_backendEn_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  payload_0_cf_pd_isRVC = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  payload_0_cf_pd_brType = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  payload_0_cf_pd_isCall = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  payload_0_cf_pd_isRet = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  payload_0_cf_pred_taken = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  payload_0_cf_storeSetHit = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  payload_0_cf_waitForRobIdx_flag = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  payload_0_cf_waitForRobIdx_value = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  payload_0_cf_loadWaitBit = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  payload_0_cf_loadWaitStrict = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  payload_0_cf_ssid = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  payload_0_cf_ftqPtr_flag = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  payload_0_cf_ftqPtr_value = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  payload_0_cf_ftqOffset = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  payload_0_ctrl_fuType = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  payload_0_ctrl_fuOpType = _RAND_18[6:0];
  _RAND_19 = {1{`RANDOM}};
  payload_0_ctrl_rfWen = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  payload_0_ctrl_fpWen = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  payload_0_ctrl_imm = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  payload_0_pdest = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  payload_0_robIdx_flag = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  payload_0_robIdx_value = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  payload_0_lqIdx_flag = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  payload_0_lqIdx_value = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  payload_0_sqIdx_flag = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  payload_0_sqIdx_value = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  payload_1_cf_foldpc = _RAND_29[9:0];
  _RAND_30 = {1{`RANDOM}};
  payload_1_cf_trigger_backendEn_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  payload_1_cf_trigger_backendEn_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  payload_1_cf_pd_isRVC = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  payload_1_cf_pd_brType = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  payload_1_cf_pd_isCall = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  payload_1_cf_pd_isRet = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  payload_1_cf_pred_taken = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  payload_1_cf_storeSetHit = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  payload_1_cf_waitForRobIdx_flag = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  payload_1_cf_waitForRobIdx_value = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  payload_1_cf_loadWaitBit = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  payload_1_cf_loadWaitStrict = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  payload_1_cf_ssid = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  payload_1_cf_ftqPtr_flag = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  payload_1_cf_ftqPtr_value = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  payload_1_cf_ftqOffset = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  payload_1_ctrl_fuType = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  payload_1_ctrl_fuOpType = _RAND_47[6:0];
  _RAND_48 = {1{`RANDOM}};
  payload_1_ctrl_rfWen = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  payload_1_ctrl_fpWen = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  payload_1_ctrl_imm = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  payload_1_pdest = _RAND_51[5:0];
  _RAND_52 = {1{`RANDOM}};
  payload_1_robIdx_flag = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  payload_1_robIdx_value = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  payload_1_lqIdx_flag = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  payload_1_lqIdx_value = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  payload_1_sqIdx_flag = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  payload_1_sqIdx_value = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  payload_2_cf_foldpc = _RAND_58[9:0];
  _RAND_59 = {1{`RANDOM}};
  payload_2_cf_trigger_backendEn_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  payload_2_cf_trigger_backendEn_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  payload_2_cf_pd_isRVC = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  payload_2_cf_pd_brType = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  payload_2_cf_pd_isCall = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  payload_2_cf_pd_isRet = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  payload_2_cf_pred_taken = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  payload_2_cf_storeSetHit = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  payload_2_cf_waitForRobIdx_flag = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  payload_2_cf_waitForRobIdx_value = _RAND_68[4:0];
  _RAND_69 = {1{`RANDOM}};
  payload_2_cf_loadWaitBit = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  payload_2_cf_loadWaitStrict = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  payload_2_cf_ssid = _RAND_71[4:0];
  _RAND_72 = {1{`RANDOM}};
  payload_2_cf_ftqPtr_flag = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  payload_2_cf_ftqPtr_value = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  payload_2_cf_ftqOffset = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  payload_2_ctrl_fuType = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  payload_2_ctrl_fuOpType = _RAND_76[6:0];
  _RAND_77 = {1{`RANDOM}};
  payload_2_ctrl_rfWen = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  payload_2_ctrl_fpWen = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  payload_2_ctrl_imm = _RAND_79[19:0];
  _RAND_80 = {1{`RANDOM}};
  payload_2_pdest = _RAND_80[5:0];
  _RAND_81 = {1{`RANDOM}};
  payload_2_robIdx_flag = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  payload_2_robIdx_value = _RAND_82[4:0];
  _RAND_83 = {1{`RANDOM}};
  payload_2_lqIdx_flag = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  payload_2_lqIdx_value = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  payload_2_sqIdx_flag = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  payload_2_sqIdx_value = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  payload_3_cf_foldpc = _RAND_87[9:0];
  _RAND_88 = {1{`RANDOM}};
  payload_3_cf_trigger_backendEn_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  payload_3_cf_trigger_backendEn_1 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  payload_3_cf_pd_isRVC = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  payload_3_cf_pd_brType = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  payload_3_cf_pd_isCall = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  payload_3_cf_pd_isRet = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  payload_3_cf_pred_taken = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  payload_3_cf_storeSetHit = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  payload_3_cf_waitForRobIdx_flag = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  payload_3_cf_waitForRobIdx_value = _RAND_97[4:0];
  _RAND_98 = {1{`RANDOM}};
  payload_3_cf_loadWaitBit = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  payload_3_cf_loadWaitStrict = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  payload_3_cf_ssid = _RAND_100[4:0];
  _RAND_101 = {1{`RANDOM}};
  payload_3_cf_ftqPtr_flag = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  payload_3_cf_ftqPtr_value = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  payload_3_cf_ftqOffset = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  payload_3_ctrl_fuType = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  payload_3_ctrl_fuOpType = _RAND_105[6:0];
  _RAND_106 = {1{`RANDOM}};
  payload_3_ctrl_rfWen = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  payload_3_ctrl_fpWen = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  payload_3_ctrl_imm = _RAND_108[19:0];
  _RAND_109 = {1{`RANDOM}};
  payload_3_pdest = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  payload_3_robIdx_flag = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  payload_3_robIdx_value = _RAND_111[4:0];
  _RAND_112 = {1{`RANDOM}};
  payload_3_lqIdx_flag = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  payload_3_lqIdx_value = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  payload_3_sqIdx_flag = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  payload_3_sqIdx_value = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  payload_4_cf_foldpc = _RAND_116[9:0];
  _RAND_117 = {1{`RANDOM}};
  payload_4_cf_trigger_backendEn_0 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  payload_4_cf_trigger_backendEn_1 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  payload_4_cf_pd_isRVC = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  payload_4_cf_pd_brType = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  payload_4_cf_pd_isCall = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  payload_4_cf_pd_isRet = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  payload_4_cf_pred_taken = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  payload_4_cf_storeSetHit = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  payload_4_cf_waitForRobIdx_flag = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  payload_4_cf_waitForRobIdx_value = _RAND_126[4:0];
  _RAND_127 = {1{`RANDOM}};
  payload_4_cf_loadWaitBit = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  payload_4_cf_loadWaitStrict = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  payload_4_cf_ssid = _RAND_129[4:0];
  _RAND_130 = {1{`RANDOM}};
  payload_4_cf_ftqPtr_flag = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  payload_4_cf_ftqPtr_value = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  payload_4_cf_ftqOffset = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  payload_4_ctrl_fuType = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  payload_4_ctrl_fuOpType = _RAND_134[6:0];
  _RAND_135 = {1{`RANDOM}};
  payload_4_ctrl_rfWen = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  payload_4_ctrl_fpWen = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  payload_4_ctrl_imm = _RAND_137[19:0];
  _RAND_138 = {1{`RANDOM}};
  payload_4_pdest = _RAND_138[5:0];
  _RAND_139 = {1{`RANDOM}};
  payload_4_robIdx_flag = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  payload_4_robIdx_value = _RAND_140[4:0];
  _RAND_141 = {1{`RANDOM}};
  payload_4_lqIdx_flag = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  payload_4_lqIdx_value = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  payload_4_sqIdx_flag = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  payload_4_sqIdx_value = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  payload_5_cf_foldpc = _RAND_145[9:0];
  _RAND_146 = {1{`RANDOM}};
  payload_5_cf_trigger_backendEn_0 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  payload_5_cf_trigger_backendEn_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  payload_5_cf_pd_isRVC = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  payload_5_cf_pd_brType = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  payload_5_cf_pd_isCall = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  payload_5_cf_pd_isRet = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  payload_5_cf_pred_taken = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  payload_5_cf_storeSetHit = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  payload_5_cf_waitForRobIdx_flag = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  payload_5_cf_waitForRobIdx_value = _RAND_155[4:0];
  _RAND_156 = {1{`RANDOM}};
  payload_5_cf_loadWaitBit = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  payload_5_cf_loadWaitStrict = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  payload_5_cf_ssid = _RAND_158[4:0];
  _RAND_159 = {1{`RANDOM}};
  payload_5_cf_ftqPtr_flag = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  payload_5_cf_ftqPtr_value = _RAND_160[2:0];
  _RAND_161 = {1{`RANDOM}};
  payload_5_cf_ftqOffset = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  payload_5_ctrl_fuType = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  payload_5_ctrl_fuOpType = _RAND_163[6:0];
  _RAND_164 = {1{`RANDOM}};
  payload_5_ctrl_rfWen = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  payload_5_ctrl_fpWen = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  payload_5_ctrl_imm = _RAND_166[19:0];
  _RAND_167 = {1{`RANDOM}};
  payload_5_pdest = _RAND_167[5:0];
  _RAND_168 = {1{`RANDOM}};
  payload_5_robIdx_flag = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  payload_5_robIdx_value = _RAND_169[4:0];
  _RAND_170 = {1{`RANDOM}};
  payload_5_lqIdx_flag = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  payload_5_lqIdx_value = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  payload_5_sqIdx_flag = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  payload_5_sqIdx_value = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  payload_6_cf_foldpc = _RAND_174[9:0];
  _RAND_175 = {1{`RANDOM}};
  payload_6_cf_trigger_backendEn_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  payload_6_cf_trigger_backendEn_1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  payload_6_cf_pd_isRVC = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  payload_6_cf_pd_brType = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  payload_6_cf_pd_isCall = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  payload_6_cf_pd_isRet = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  payload_6_cf_pred_taken = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  payload_6_cf_storeSetHit = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  payload_6_cf_waitForRobIdx_flag = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  payload_6_cf_waitForRobIdx_value = _RAND_184[4:0];
  _RAND_185 = {1{`RANDOM}};
  payload_6_cf_loadWaitBit = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  payload_6_cf_loadWaitStrict = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  payload_6_cf_ssid = _RAND_187[4:0];
  _RAND_188 = {1{`RANDOM}};
  payload_6_cf_ftqPtr_flag = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  payload_6_cf_ftqPtr_value = _RAND_189[2:0];
  _RAND_190 = {1{`RANDOM}};
  payload_6_cf_ftqOffset = _RAND_190[2:0];
  _RAND_191 = {1{`RANDOM}};
  payload_6_ctrl_fuType = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  payload_6_ctrl_fuOpType = _RAND_192[6:0];
  _RAND_193 = {1{`RANDOM}};
  payload_6_ctrl_rfWen = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  payload_6_ctrl_fpWen = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  payload_6_ctrl_imm = _RAND_195[19:0];
  _RAND_196 = {1{`RANDOM}};
  payload_6_pdest = _RAND_196[5:0];
  _RAND_197 = {1{`RANDOM}};
  payload_6_robIdx_flag = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  payload_6_robIdx_value = _RAND_198[4:0];
  _RAND_199 = {1{`RANDOM}};
  payload_6_lqIdx_flag = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  payload_6_lqIdx_value = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  payload_6_sqIdx_flag = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  payload_6_sqIdx_value = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  payload_7_cf_foldpc = _RAND_203[9:0];
  _RAND_204 = {1{`RANDOM}};
  payload_7_cf_trigger_backendEn_0 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  payload_7_cf_trigger_backendEn_1 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  payload_7_cf_pd_isRVC = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  payload_7_cf_pd_brType = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  payload_7_cf_pd_isCall = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  payload_7_cf_pd_isRet = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  payload_7_cf_pred_taken = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  payload_7_cf_storeSetHit = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  payload_7_cf_waitForRobIdx_flag = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  payload_7_cf_waitForRobIdx_value = _RAND_213[4:0];
  _RAND_214 = {1{`RANDOM}};
  payload_7_cf_loadWaitBit = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  payload_7_cf_loadWaitStrict = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  payload_7_cf_ssid = _RAND_216[4:0];
  _RAND_217 = {1{`RANDOM}};
  payload_7_cf_ftqPtr_flag = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  payload_7_cf_ftqPtr_value = _RAND_218[2:0];
  _RAND_219 = {1{`RANDOM}};
  payload_7_cf_ftqOffset = _RAND_219[2:0];
  _RAND_220 = {1{`RANDOM}};
  payload_7_ctrl_fuType = _RAND_220[3:0];
  _RAND_221 = {1{`RANDOM}};
  payload_7_ctrl_fuOpType = _RAND_221[6:0];
  _RAND_222 = {1{`RANDOM}};
  payload_7_ctrl_rfWen = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  payload_7_ctrl_fpWen = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  payload_7_ctrl_imm = _RAND_224[19:0];
  _RAND_225 = {1{`RANDOM}};
  payload_7_pdest = _RAND_225[5:0];
  _RAND_226 = {1{`RANDOM}};
  payload_7_robIdx_flag = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  payload_7_robIdx_value = _RAND_227[4:0];
  _RAND_228 = {1{`RANDOM}};
  payload_7_lqIdx_flag = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  payload_7_lqIdx_value = _RAND_229[3:0];
  _RAND_230 = {1{`RANDOM}};
  payload_7_sqIdx_flag = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  payload_7_sqIdx_value = _RAND_231[3:0];
  _RAND_232 = {1{`RANDOM}};
  payload_8_cf_foldpc = _RAND_232[9:0];
  _RAND_233 = {1{`RANDOM}};
  payload_8_cf_trigger_backendEn_0 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  payload_8_cf_trigger_backendEn_1 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  payload_8_cf_pd_isRVC = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  payload_8_cf_pd_brType = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  payload_8_cf_pd_isCall = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  payload_8_cf_pd_isRet = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  payload_8_cf_pred_taken = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  payload_8_cf_storeSetHit = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  payload_8_cf_waitForRobIdx_flag = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  payload_8_cf_waitForRobIdx_value = _RAND_242[4:0];
  _RAND_243 = {1{`RANDOM}};
  payload_8_cf_loadWaitBit = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  payload_8_cf_loadWaitStrict = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  payload_8_cf_ssid = _RAND_245[4:0];
  _RAND_246 = {1{`RANDOM}};
  payload_8_cf_ftqPtr_flag = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  payload_8_cf_ftqPtr_value = _RAND_247[2:0];
  _RAND_248 = {1{`RANDOM}};
  payload_8_cf_ftqOffset = _RAND_248[2:0];
  _RAND_249 = {1{`RANDOM}};
  payload_8_ctrl_fuType = _RAND_249[3:0];
  _RAND_250 = {1{`RANDOM}};
  payload_8_ctrl_fuOpType = _RAND_250[6:0];
  _RAND_251 = {1{`RANDOM}};
  payload_8_ctrl_rfWen = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  payload_8_ctrl_fpWen = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  payload_8_ctrl_imm = _RAND_253[19:0];
  _RAND_254 = {1{`RANDOM}};
  payload_8_pdest = _RAND_254[5:0];
  _RAND_255 = {1{`RANDOM}};
  payload_8_robIdx_flag = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  payload_8_robIdx_value = _RAND_256[4:0];
  _RAND_257 = {1{`RANDOM}};
  payload_8_lqIdx_flag = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  payload_8_lqIdx_value = _RAND_258[3:0];
  _RAND_259 = {1{`RANDOM}};
  payload_8_sqIdx_flag = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  payload_8_sqIdx_value = _RAND_260[3:0];
  _RAND_261 = {1{`RANDOM}};
  payload_9_cf_foldpc = _RAND_261[9:0];
  _RAND_262 = {1{`RANDOM}};
  payload_9_cf_trigger_backendEn_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  payload_9_cf_trigger_backendEn_1 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  payload_9_cf_pd_isRVC = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  payload_9_cf_pd_brType = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  payload_9_cf_pd_isCall = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  payload_9_cf_pd_isRet = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  payload_9_cf_pred_taken = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  payload_9_cf_storeSetHit = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  payload_9_cf_waitForRobIdx_flag = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  payload_9_cf_waitForRobIdx_value = _RAND_271[4:0];
  _RAND_272 = {1{`RANDOM}};
  payload_9_cf_loadWaitBit = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  payload_9_cf_loadWaitStrict = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  payload_9_cf_ssid = _RAND_274[4:0];
  _RAND_275 = {1{`RANDOM}};
  payload_9_cf_ftqPtr_flag = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  payload_9_cf_ftqPtr_value = _RAND_276[2:0];
  _RAND_277 = {1{`RANDOM}};
  payload_9_cf_ftqOffset = _RAND_277[2:0];
  _RAND_278 = {1{`RANDOM}};
  payload_9_ctrl_fuType = _RAND_278[3:0];
  _RAND_279 = {1{`RANDOM}};
  payload_9_ctrl_fuOpType = _RAND_279[6:0];
  _RAND_280 = {1{`RANDOM}};
  payload_9_ctrl_rfWen = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  payload_9_ctrl_fpWen = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  payload_9_ctrl_imm = _RAND_282[19:0];
  _RAND_283 = {1{`RANDOM}};
  payload_9_pdest = _RAND_283[5:0];
  _RAND_284 = {1{`RANDOM}};
  payload_9_robIdx_flag = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  payload_9_robIdx_value = _RAND_285[4:0];
  _RAND_286 = {1{`RANDOM}};
  payload_9_lqIdx_flag = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  payload_9_lqIdx_value = _RAND_287[3:0];
  _RAND_288 = {1{`RANDOM}};
  payload_9_sqIdx_flag = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  payload_9_sqIdx_value = _RAND_289[3:0];
  _RAND_290 = {1{`RANDOM}};
  payload_10_cf_foldpc = _RAND_290[9:0];
  _RAND_291 = {1{`RANDOM}};
  payload_10_cf_trigger_backendEn_0 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  payload_10_cf_trigger_backendEn_1 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  payload_10_cf_pd_isRVC = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  payload_10_cf_pd_brType = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  payload_10_cf_pd_isCall = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  payload_10_cf_pd_isRet = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  payload_10_cf_pred_taken = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  payload_10_cf_storeSetHit = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  payload_10_cf_waitForRobIdx_flag = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  payload_10_cf_waitForRobIdx_value = _RAND_300[4:0];
  _RAND_301 = {1{`RANDOM}};
  payload_10_cf_loadWaitBit = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  payload_10_cf_loadWaitStrict = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  payload_10_cf_ssid = _RAND_303[4:0];
  _RAND_304 = {1{`RANDOM}};
  payload_10_cf_ftqPtr_flag = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  payload_10_cf_ftqPtr_value = _RAND_305[2:0];
  _RAND_306 = {1{`RANDOM}};
  payload_10_cf_ftqOffset = _RAND_306[2:0];
  _RAND_307 = {1{`RANDOM}};
  payload_10_ctrl_fuType = _RAND_307[3:0];
  _RAND_308 = {1{`RANDOM}};
  payload_10_ctrl_fuOpType = _RAND_308[6:0];
  _RAND_309 = {1{`RANDOM}};
  payload_10_ctrl_rfWen = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  payload_10_ctrl_fpWen = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  payload_10_ctrl_imm = _RAND_311[19:0];
  _RAND_312 = {1{`RANDOM}};
  payload_10_pdest = _RAND_312[5:0];
  _RAND_313 = {1{`RANDOM}};
  payload_10_robIdx_flag = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  payload_10_robIdx_value = _RAND_314[4:0];
  _RAND_315 = {1{`RANDOM}};
  payload_10_lqIdx_flag = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  payload_10_lqIdx_value = _RAND_316[3:0];
  _RAND_317 = {1{`RANDOM}};
  payload_10_sqIdx_flag = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  payload_10_sqIdx_value = _RAND_318[3:0];
  _RAND_319 = {1{`RANDOM}};
  payload_11_cf_foldpc = _RAND_319[9:0];
  _RAND_320 = {1{`RANDOM}};
  payload_11_cf_trigger_backendEn_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  payload_11_cf_trigger_backendEn_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  payload_11_cf_pd_isRVC = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  payload_11_cf_pd_brType = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  payload_11_cf_pd_isCall = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  payload_11_cf_pd_isRet = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  payload_11_cf_pred_taken = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  payload_11_cf_storeSetHit = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  payload_11_cf_waitForRobIdx_flag = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  payload_11_cf_waitForRobIdx_value = _RAND_329[4:0];
  _RAND_330 = {1{`RANDOM}};
  payload_11_cf_loadWaitBit = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  payload_11_cf_loadWaitStrict = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  payload_11_cf_ssid = _RAND_332[4:0];
  _RAND_333 = {1{`RANDOM}};
  payload_11_cf_ftqPtr_flag = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  payload_11_cf_ftqPtr_value = _RAND_334[2:0];
  _RAND_335 = {1{`RANDOM}};
  payload_11_cf_ftqOffset = _RAND_335[2:0];
  _RAND_336 = {1{`RANDOM}};
  payload_11_ctrl_fuType = _RAND_336[3:0];
  _RAND_337 = {1{`RANDOM}};
  payload_11_ctrl_fuOpType = _RAND_337[6:0];
  _RAND_338 = {1{`RANDOM}};
  payload_11_ctrl_rfWen = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  payload_11_ctrl_fpWen = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  payload_11_ctrl_imm = _RAND_340[19:0];
  _RAND_341 = {1{`RANDOM}};
  payload_11_pdest = _RAND_341[5:0];
  _RAND_342 = {1{`RANDOM}};
  payload_11_robIdx_flag = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  payload_11_robIdx_value = _RAND_343[4:0];
  _RAND_344 = {1{`RANDOM}};
  payload_11_lqIdx_flag = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  payload_11_lqIdx_value = _RAND_345[3:0];
  _RAND_346 = {1{`RANDOM}};
  payload_11_sqIdx_flag = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  payload_11_sqIdx_value = _RAND_347[3:0];
  _RAND_348 = {1{`RANDOM}};
  payload_12_cf_foldpc = _RAND_348[9:0];
  _RAND_349 = {1{`RANDOM}};
  payload_12_cf_trigger_backendEn_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  payload_12_cf_trigger_backendEn_1 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  payload_12_cf_pd_isRVC = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  payload_12_cf_pd_brType = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  payload_12_cf_pd_isCall = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  payload_12_cf_pd_isRet = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  payload_12_cf_pred_taken = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  payload_12_cf_storeSetHit = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  payload_12_cf_waitForRobIdx_flag = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  payload_12_cf_waitForRobIdx_value = _RAND_358[4:0];
  _RAND_359 = {1{`RANDOM}};
  payload_12_cf_loadWaitBit = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  payload_12_cf_loadWaitStrict = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  payload_12_cf_ssid = _RAND_361[4:0];
  _RAND_362 = {1{`RANDOM}};
  payload_12_cf_ftqPtr_flag = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  payload_12_cf_ftqPtr_value = _RAND_363[2:0];
  _RAND_364 = {1{`RANDOM}};
  payload_12_cf_ftqOffset = _RAND_364[2:0];
  _RAND_365 = {1{`RANDOM}};
  payload_12_ctrl_fuType = _RAND_365[3:0];
  _RAND_366 = {1{`RANDOM}};
  payload_12_ctrl_fuOpType = _RAND_366[6:0];
  _RAND_367 = {1{`RANDOM}};
  payload_12_ctrl_rfWen = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  payload_12_ctrl_fpWen = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  payload_12_ctrl_imm = _RAND_369[19:0];
  _RAND_370 = {1{`RANDOM}};
  payload_12_pdest = _RAND_370[5:0];
  _RAND_371 = {1{`RANDOM}};
  payload_12_robIdx_flag = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  payload_12_robIdx_value = _RAND_372[4:0];
  _RAND_373 = {1{`RANDOM}};
  payload_12_lqIdx_flag = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  payload_12_lqIdx_value = _RAND_374[3:0];
  _RAND_375 = {1{`RANDOM}};
  payload_12_sqIdx_flag = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  payload_12_sqIdx_value = _RAND_376[3:0];
  _RAND_377 = {1{`RANDOM}};
  payload_13_cf_foldpc = _RAND_377[9:0];
  _RAND_378 = {1{`RANDOM}};
  payload_13_cf_trigger_backendEn_0 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  payload_13_cf_trigger_backendEn_1 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  payload_13_cf_pd_isRVC = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  payload_13_cf_pd_brType = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  payload_13_cf_pd_isCall = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  payload_13_cf_pd_isRet = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  payload_13_cf_pred_taken = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  payload_13_cf_storeSetHit = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  payload_13_cf_waitForRobIdx_flag = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  payload_13_cf_waitForRobIdx_value = _RAND_387[4:0];
  _RAND_388 = {1{`RANDOM}};
  payload_13_cf_loadWaitBit = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  payload_13_cf_loadWaitStrict = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  payload_13_cf_ssid = _RAND_390[4:0];
  _RAND_391 = {1{`RANDOM}};
  payload_13_cf_ftqPtr_flag = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  payload_13_cf_ftqPtr_value = _RAND_392[2:0];
  _RAND_393 = {1{`RANDOM}};
  payload_13_cf_ftqOffset = _RAND_393[2:0];
  _RAND_394 = {1{`RANDOM}};
  payload_13_ctrl_fuType = _RAND_394[3:0];
  _RAND_395 = {1{`RANDOM}};
  payload_13_ctrl_fuOpType = _RAND_395[6:0];
  _RAND_396 = {1{`RANDOM}};
  payload_13_ctrl_rfWen = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  payload_13_ctrl_fpWen = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  payload_13_ctrl_imm = _RAND_398[19:0];
  _RAND_399 = {1{`RANDOM}};
  payload_13_pdest = _RAND_399[5:0];
  _RAND_400 = {1{`RANDOM}};
  payload_13_robIdx_flag = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  payload_13_robIdx_value = _RAND_401[4:0];
  _RAND_402 = {1{`RANDOM}};
  payload_13_lqIdx_flag = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  payload_13_lqIdx_value = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  payload_13_sqIdx_flag = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  payload_13_sqIdx_value = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  payload_14_cf_foldpc = _RAND_406[9:0];
  _RAND_407 = {1{`RANDOM}};
  payload_14_cf_trigger_backendEn_0 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  payload_14_cf_trigger_backendEn_1 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  payload_14_cf_pd_isRVC = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  payload_14_cf_pd_brType = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  payload_14_cf_pd_isCall = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  payload_14_cf_pd_isRet = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  payload_14_cf_pred_taken = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  payload_14_cf_storeSetHit = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  payload_14_cf_waitForRobIdx_flag = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  payload_14_cf_waitForRobIdx_value = _RAND_416[4:0];
  _RAND_417 = {1{`RANDOM}};
  payload_14_cf_loadWaitBit = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  payload_14_cf_loadWaitStrict = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  payload_14_cf_ssid = _RAND_419[4:0];
  _RAND_420 = {1{`RANDOM}};
  payload_14_cf_ftqPtr_flag = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  payload_14_cf_ftqPtr_value = _RAND_421[2:0];
  _RAND_422 = {1{`RANDOM}};
  payload_14_cf_ftqOffset = _RAND_422[2:0];
  _RAND_423 = {1{`RANDOM}};
  payload_14_ctrl_fuType = _RAND_423[3:0];
  _RAND_424 = {1{`RANDOM}};
  payload_14_ctrl_fuOpType = _RAND_424[6:0];
  _RAND_425 = {1{`RANDOM}};
  payload_14_ctrl_rfWen = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  payload_14_ctrl_fpWen = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  payload_14_ctrl_imm = _RAND_427[19:0];
  _RAND_428 = {1{`RANDOM}};
  payload_14_pdest = _RAND_428[5:0];
  _RAND_429 = {1{`RANDOM}};
  payload_14_robIdx_flag = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  payload_14_robIdx_value = _RAND_430[4:0];
  _RAND_431 = {1{`RANDOM}};
  payload_14_lqIdx_flag = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  payload_14_lqIdx_value = _RAND_432[3:0];
  _RAND_433 = {1{`RANDOM}};
  payload_14_sqIdx_flag = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  payload_14_sqIdx_value = _RAND_434[3:0];
  _RAND_435 = {1{`RANDOM}};
  payload_15_cf_foldpc = _RAND_435[9:0];
  _RAND_436 = {1{`RANDOM}};
  payload_15_cf_trigger_backendEn_0 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  payload_15_cf_trigger_backendEn_1 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  payload_15_cf_pd_isRVC = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  payload_15_cf_pd_brType = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  payload_15_cf_pd_isCall = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  payload_15_cf_pd_isRet = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  payload_15_cf_pred_taken = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  payload_15_cf_storeSetHit = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  payload_15_cf_waitForRobIdx_flag = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  payload_15_cf_waitForRobIdx_value = _RAND_445[4:0];
  _RAND_446 = {1{`RANDOM}};
  payload_15_cf_loadWaitBit = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  payload_15_cf_loadWaitStrict = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  payload_15_cf_ssid = _RAND_448[4:0];
  _RAND_449 = {1{`RANDOM}};
  payload_15_cf_ftqPtr_flag = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  payload_15_cf_ftqPtr_value = _RAND_450[2:0];
  _RAND_451 = {1{`RANDOM}};
  payload_15_cf_ftqOffset = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  payload_15_ctrl_fuType = _RAND_452[3:0];
  _RAND_453 = {1{`RANDOM}};
  payload_15_ctrl_fuOpType = _RAND_453[6:0];
  _RAND_454 = {1{`RANDOM}};
  payload_15_ctrl_rfWen = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  payload_15_ctrl_fpWen = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  payload_15_ctrl_imm = _RAND_456[19:0];
  _RAND_457 = {1{`RANDOM}};
  payload_15_pdest = _RAND_457[5:0];
  _RAND_458 = {1{`RANDOM}};
  payload_15_robIdx_flag = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  payload_15_robIdx_value = _RAND_459[4:0];
  _RAND_460 = {1{`RANDOM}};
  payload_15_lqIdx_flag = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  payload_15_lqIdx_value = _RAND_461[3:0];
  _RAND_462 = {1{`RANDOM}};
  payload_15_sqIdx_flag = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  payload_15_sqIdx_value = _RAND_463[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

