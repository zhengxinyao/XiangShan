module SbufferData(
  input          clock,
  input          reset,
  input          io_writeReq_0_valid,
  input  [3:0]   io_writeReq_0_bits_wvec,
  input  [15:0]  io_writeReq_0_bits_mask,
  input  [127:0] io_writeReq_0_bits_data,
  input  [31:0]  io_writeReq_0_bits_vwordOffset,
  input          io_writeReq_0_bits_wline,
  input          io_writeReq_1_valid,
  input  [3:0]   io_writeReq_1_bits_wvec,
  input  [15:0]  io_writeReq_1_bits_mask,
  input  [127:0] io_writeReq_1_bits_data,
  input  [31:0]  io_writeReq_1_bits_vwordOffset,
  input          io_writeReq_1_bits_wline,
  input          io_maskFlushReq_0_valid,
  input  [3:0]   io_maskFlushReq_0_bits_wvec,
  input          io_maskFlushReq_1_valid,
  input  [3:0]   io_maskFlushReq_1_bits_wvec,
  output [7:0]   io_dataOut_0_0_0,
  output [7:0]   io_dataOut_0_0_1,
  output [7:0]   io_dataOut_0_0_2,
  output [7:0]   io_dataOut_0_0_3,
  output [7:0]   io_dataOut_0_0_4,
  output [7:0]   io_dataOut_0_0_5,
  output [7:0]   io_dataOut_0_0_6,
  output [7:0]   io_dataOut_0_0_7,
  output [7:0]   io_dataOut_0_0_8,
  output [7:0]   io_dataOut_0_0_9,
  output [7:0]   io_dataOut_0_0_10,
  output [7:0]   io_dataOut_0_0_11,
  output [7:0]   io_dataOut_0_0_12,
  output [7:0]   io_dataOut_0_0_13,
  output [7:0]   io_dataOut_0_0_14,
  output [7:0]   io_dataOut_0_0_15,
  output [7:0]   io_dataOut_0_1_0,
  output [7:0]   io_dataOut_0_1_1,
  output [7:0]   io_dataOut_0_1_2,
  output [7:0]   io_dataOut_0_1_3,
  output [7:0]   io_dataOut_0_1_4,
  output [7:0]   io_dataOut_0_1_5,
  output [7:0]   io_dataOut_0_1_6,
  output [7:0]   io_dataOut_0_1_7,
  output [7:0]   io_dataOut_0_1_8,
  output [7:0]   io_dataOut_0_1_9,
  output [7:0]   io_dataOut_0_1_10,
  output [7:0]   io_dataOut_0_1_11,
  output [7:0]   io_dataOut_0_1_12,
  output [7:0]   io_dataOut_0_1_13,
  output [7:0]   io_dataOut_0_1_14,
  output [7:0]   io_dataOut_0_1_15,
  output [7:0]   io_dataOut_0_2_0,
  output [7:0]   io_dataOut_0_2_1,
  output [7:0]   io_dataOut_0_2_2,
  output [7:0]   io_dataOut_0_2_3,
  output [7:0]   io_dataOut_0_2_4,
  output [7:0]   io_dataOut_0_2_5,
  output [7:0]   io_dataOut_0_2_6,
  output [7:0]   io_dataOut_0_2_7,
  output [7:0]   io_dataOut_0_2_8,
  output [7:0]   io_dataOut_0_2_9,
  output [7:0]   io_dataOut_0_2_10,
  output [7:0]   io_dataOut_0_2_11,
  output [7:0]   io_dataOut_0_2_12,
  output [7:0]   io_dataOut_0_2_13,
  output [7:0]   io_dataOut_0_2_14,
  output [7:0]   io_dataOut_0_2_15,
  output [7:0]   io_dataOut_0_3_0,
  output [7:0]   io_dataOut_0_3_1,
  output [7:0]   io_dataOut_0_3_2,
  output [7:0]   io_dataOut_0_3_3,
  output [7:0]   io_dataOut_0_3_4,
  output [7:0]   io_dataOut_0_3_5,
  output [7:0]   io_dataOut_0_3_6,
  output [7:0]   io_dataOut_0_3_7,
  output [7:0]   io_dataOut_0_3_8,
  output [7:0]   io_dataOut_0_3_9,
  output [7:0]   io_dataOut_0_3_10,
  output [7:0]   io_dataOut_0_3_11,
  output [7:0]   io_dataOut_0_3_12,
  output [7:0]   io_dataOut_0_3_13,
  output [7:0]   io_dataOut_0_3_14,
  output [7:0]   io_dataOut_0_3_15,
  output [7:0]   io_dataOut_1_0_0,
  output [7:0]   io_dataOut_1_0_1,
  output [7:0]   io_dataOut_1_0_2,
  output [7:0]   io_dataOut_1_0_3,
  output [7:0]   io_dataOut_1_0_4,
  output [7:0]   io_dataOut_1_0_5,
  output [7:0]   io_dataOut_1_0_6,
  output [7:0]   io_dataOut_1_0_7,
  output [7:0]   io_dataOut_1_0_8,
  output [7:0]   io_dataOut_1_0_9,
  output [7:0]   io_dataOut_1_0_10,
  output [7:0]   io_dataOut_1_0_11,
  output [7:0]   io_dataOut_1_0_12,
  output [7:0]   io_dataOut_1_0_13,
  output [7:0]   io_dataOut_1_0_14,
  output [7:0]   io_dataOut_1_0_15,
  output [7:0]   io_dataOut_1_1_0,
  output [7:0]   io_dataOut_1_1_1,
  output [7:0]   io_dataOut_1_1_2,
  output [7:0]   io_dataOut_1_1_3,
  output [7:0]   io_dataOut_1_1_4,
  output [7:0]   io_dataOut_1_1_5,
  output [7:0]   io_dataOut_1_1_6,
  output [7:0]   io_dataOut_1_1_7,
  output [7:0]   io_dataOut_1_1_8,
  output [7:0]   io_dataOut_1_1_9,
  output [7:0]   io_dataOut_1_1_10,
  output [7:0]   io_dataOut_1_1_11,
  output [7:0]   io_dataOut_1_1_12,
  output [7:0]   io_dataOut_1_1_13,
  output [7:0]   io_dataOut_1_1_14,
  output [7:0]   io_dataOut_1_1_15,
  output [7:0]   io_dataOut_1_2_0,
  output [7:0]   io_dataOut_1_2_1,
  output [7:0]   io_dataOut_1_2_2,
  output [7:0]   io_dataOut_1_2_3,
  output [7:0]   io_dataOut_1_2_4,
  output [7:0]   io_dataOut_1_2_5,
  output [7:0]   io_dataOut_1_2_6,
  output [7:0]   io_dataOut_1_2_7,
  output [7:0]   io_dataOut_1_2_8,
  output [7:0]   io_dataOut_1_2_9,
  output [7:0]   io_dataOut_1_2_10,
  output [7:0]   io_dataOut_1_2_11,
  output [7:0]   io_dataOut_1_2_12,
  output [7:0]   io_dataOut_1_2_13,
  output [7:0]   io_dataOut_1_2_14,
  output [7:0]   io_dataOut_1_2_15,
  output [7:0]   io_dataOut_1_3_0,
  output [7:0]   io_dataOut_1_3_1,
  output [7:0]   io_dataOut_1_3_2,
  output [7:0]   io_dataOut_1_3_3,
  output [7:0]   io_dataOut_1_3_4,
  output [7:0]   io_dataOut_1_3_5,
  output [7:0]   io_dataOut_1_3_6,
  output [7:0]   io_dataOut_1_3_7,
  output [7:0]   io_dataOut_1_3_8,
  output [7:0]   io_dataOut_1_3_9,
  output [7:0]   io_dataOut_1_3_10,
  output [7:0]   io_dataOut_1_3_11,
  output [7:0]   io_dataOut_1_3_12,
  output [7:0]   io_dataOut_1_3_13,
  output [7:0]   io_dataOut_1_3_14,
  output [7:0]   io_dataOut_1_3_15,
  output [7:0]   io_dataOut_2_0_0,
  output [7:0]   io_dataOut_2_0_1,
  output [7:0]   io_dataOut_2_0_2,
  output [7:0]   io_dataOut_2_0_3,
  output [7:0]   io_dataOut_2_0_4,
  output [7:0]   io_dataOut_2_0_5,
  output [7:0]   io_dataOut_2_0_6,
  output [7:0]   io_dataOut_2_0_7,
  output [7:0]   io_dataOut_2_0_8,
  output [7:0]   io_dataOut_2_0_9,
  output [7:0]   io_dataOut_2_0_10,
  output [7:0]   io_dataOut_2_0_11,
  output [7:0]   io_dataOut_2_0_12,
  output [7:0]   io_dataOut_2_0_13,
  output [7:0]   io_dataOut_2_0_14,
  output [7:0]   io_dataOut_2_0_15,
  output [7:0]   io_dataOut_2_1_0,
  output [7:0]   io_dataOut_2_1_1,
  output [7:0]   io_dataOut_2_1_2,
  output [7:0]   io_dataOut_2_1_3,
  output [7:0]   io_dataOut_2_1_4,
  output [7:0]   io_dataOut_2_1_5,
  output [7:0]   io_dataOut_2_1_6,
  output [7:0]   io_dataOut_2_1_7,
  output [7:0]   io_dataOut_2_1_8,
  output [7:0]   io_dataOut_2_1_9,
  output [7:0]   io_dataOut_2_1_10,
  output [7:0]   io_dataOut_2_1_11,
  output [7:0]   io_dataOut_2_1_12,
  output [7:0]   io_dataOut_2_1_13,
  output [7:0]   io_dataOut_2_1_14,
  output [7:0]   io_dataOut_2_1_15,
  output [7:0]   io_dataOut_2_2_0,
  output [7:0]   io_dataOut_2_2_1,
  output [7:0]   io_dataOut_2_2_2,
  output [7:0]   io_dataOut_2_2_3,
  output [7:0]   io_dataOut_2_2_4,
  output [7:0]   io_dataOut_2_2_5,
  output [7:0]   io_dataOut_2_2_6,
  output [7:0]   io_dataOut_2_2_7,
  output [7:0]   io_dataOut_2_2_8,
  output [7:0]   io_dataOut_2_2_9,
  output [7:0]   io_dataOut_2_2_10,
  output [7:0]   io_dataOut_2_2_11,
  output [7:0]   io_dataOut_2_2_12,
  output [7:0]   io_dataOut_2_2_13,
  output [7:0]   io_dataOut_2_2_14,
  output [7:0]   io_dataOut_2_2_15,
  output [7:0]   io_dataOut_2_3_0,
  output [7:0]   io_dataOut_2_3_1,
  output [7:0]   io_dataOut_2_3_2,
  output [7:0]   io_dataOut_2_3_3,
  output [7:0]   io_dataOut_2_3_4,
  output [7:0]   io_dataOut_2_3_5,
  output [7:0]   io_dataOut_2_3_6,
  output [7:0]   io_dataOut_2_3_7,
  output [7:0]   io_dataOut_2_3_8,
  output [7:0]   io_dataOut_2_3_9,
  output [7:0]   io_dataOut_2_3_10,
  output [7:0]   io_dataOut_2_3_11,
  output [7:0]   io_dataOut_2_3_12,
  output [7:0]   io_dataOut_2_3_13,
  output [7:0]   io_dataOut_2_3_14,
  output [7:0]   io_dataOut_2_3_15,
  output [7:0]   io_dataOut_3_0_0,
  output [7:0]   io_dataOut_3_0_1,
  output [7:0]   io_dataOut_3_0_2,
  output [7:0]   io_dataOut_3_0_3,
  output [7:0]   io_dataOut_3_0_4,
  output [7:0]   io_dataOut_3_0_5,
  output [7:0]   io_dataOut_3_0_6,
  output [7:0]   io_dataOut_3_0_7,
  output [7:0]   io_dataOut_3_0_8,
  output [7:0]   io_dataOut_3_0_9,
  output [7:0]   io_dataOut_3_0_10,
  output [7:0]   io_dataOut_3_0_11,
  output [7:0]   io_dataOut_3_0_12,
  output [7:0]   io_dataOut_3_0_13,
  output [7:0]   io_dataOut_3_0_14,
  output [7:0]   io_dataOut_3_0_15,
  output [7:0]   io_dataOut_3_1_0,
  output [7:0]   io_dataOut_3_1_1,
  output [7:0]   io_dataOut_3_1_2,
  output [7:0]   io_dataOut_3_1_3,
  output [7:0]   io_dataOut_3_1_4,
  output [7:0]   io_dataOut_3_1_5,
  output [7:0]   io_dataOut_3_1_6,
  output [7:0]   io_dataOut_3_1_7,
  output [7:0]   io_dataOut_3_1_8,
  output [7:0]   io_dataOut_3_1_9,
  output [7:0]   io_dataOut_3_1_10,
  output [7:0]   io_dataOut_3_1_11,
  output [7:0]   io_dataOut_3_1_12,
  output [7:0]   io_dataOut_3_1_13,
  output [7:0]   io_dataOut_3_1_14,
  output [7:0]   io_dataOut_3_1_15,
  output [7:0]   io_dataOut_3_2_0,
  output [7:0]   io_dataOut_3_2_1,
  output [7:0]   io_dataOut_3_2_2,
  output [7:0]   io_dataOut_3_2_3,
  output [7:0]   io_dataOut_3_2_4,
  output [7:0]   io_dataOut_3_2_5,
  output [7:0]   io_dataOut_3_2_6,
  output [7:0]   io_dataOut_3_2_7,
  output [7:0]   io_dataOut_3_2_8,
  output [7:0]   io_dataOut_3_2_9,
  output [7:0]   io_dataOut_3_2_10,
  output [7:0]   io_dataOut_3_2_11,
  output [7:0]   io_dataOut_3_2_12,
  output [7:0]   io_dataOut_3_2_13,
  output [7:0]   io_dataOut_3_2_14,
  output [7:0]   io_dataOut_3_2_15,
  output [7:0]   io_dataOut_3_3_0,
  output [7:0]   io_dataOut_3_3_1,
  output [7:0]   io_dataOut_3_3_2,
  output [7:0]   io_dataOut_3_3_3,
  output [7:0]   io_dataOut_3_3_4,
  output [7:0]   io_dataOut_3_3_5,
  output [7:0]   io_dataOut_3_3_6,
  output [7:0]   io_dataOut_3_3_7,
  output [7:0]   io_dataOut_3_3_8,
  output [7:0]   io_dataOut_3_3_9,
  output [7:0]   io_dataOut_3_3_10,
  output [7:0]   io_dataOut_3_3_11,
  output [7:0]   io_dataOut_3_3_12,
  output [7:0]   io_dataOut_3_3_13,
  output [7:0]   io_dataOut_3_3_14,
  output [7:0]   io_dataOut_3_3_15,
  output         io_maskOut_0_0_0,
  output         io_maskOut_0_0_1,
  output         io_maskOut_0_0_2,
  output         io_maskOut_0_0_3,
  output         io_maskOut_0_0_4,
  output         io_maskOut_0_0_5,
  output         io_maskOut_0_0_6,
  output         io_maskOut_0_0_7,
  output         io_maskOut_0_0_8,
  output         io_maskOut_0_0_9,
  output         io_maskOut_0_0_10,
  output         io_maskOut_0_0_11,
  output         io_maskOut_0_0_12,
  output         io_maskOut_0_0_13,
  output         io_maskOut_0_0_14,
  output         io_maskOut_0_0_15,
  output         io_maskOut_0_1_0,
  output         io_maskOut_0_1_1,
  output         io_maskOut_0_1_2,
  output         io_maskOut_0_1_3,
  output         io_maskOut_0_1_4,
  output         io_maskOut_0_1_5,
  output         io_maskOut_0_1_6,
  output         io_maskOut_0_1_7,
  output         io_maskOut_0_1_8,
  output         io_maskOut_0_1_9,
  output         io_maskOut_0_1_10,
  output         io_maskOut_0_1_11,
  output         io_maskOut_0_1_12,
  output         io_maskOut_0_1_13,
  output         io_maskOut_0_1_14,
  output         io_maskOut_0_1_15,
  output         io_maskOut_0_2_0,
  output         io_maskOut_0_2_1,
  output         io_maskOut_0_2_2,
  output         io_maskOut_0_2_3,
  output         io_maskOut_0_2_4,
  output         io_maskOut_0_2_5,
  output         io_maskOut_0_2_6,
  output         io_maskOut_0_2_7,
  output         io_maskOut_0_2_8,
  output         io_maskOut_0_2_9,
  output         io_maskOut_0_2_10,
  output         io_maskOut_0_2_11,
  output         io_maskOut_0_2_12,
  output         io_maskOut_0_2_13,
  output         io_maskOut_0_2_14,
  output         io_maskOut_0_2_15,
  output         io_maskOut_0_3_0,
  output         io_maskOut_0_3_1,
  output         io_maskOut_0_3_2,
  output         io_maskOut_0_3_3,
  output         io_maskOut_0_3_4,
  output         io_maskOut_0_3_5,
  output         io_maskOut_0_3_6,
  output         io_maskOut_0_3_7,
  output         io_maskOut_0_3_8,
  output         io_maskOut_0_3_9,
  output         io_maskOut_0_3_10,
  output         io_maskOut_0_3_11,
  output         io_maskOut_0_3_12,
  output         io_maskOut_0_3_13,
  output         io_maskOut_0_3_14,
  output         io_maskOut_0_3_15,
  output         io_maskOut_1_0_0,
  output         io_maskOut_1_0_1,
  output         io_maskOut_1_0_2,
  output         io_maskOut_1_0_3,
  output         io_maskOut_1_0_4,
  output         io_maskOut_1_0_5,
  output         io_maskOut_1_0_6,
  output         io_maskOut_1_0_7,
  output         io_maskOut_1_0_8,
  output         io_maskOut_1_0_9,
  output         io_maskOut_1_0_10,
  output         io_maskOut_1_0_11,
  output         io_maskOut_1_0_12,
  output         io_maskOut_1_0_13,
  output         io_maskOut_1_0_14,
  output         io_maskOut_1_0_15,
  output         io_maskOut_1_1_0,
  output         io_maskOut_1_1_1,
  output         io_maskOut_1_1_2,
  output         io_maskOut_1_1_3,
  output         io_maskOut_1_1_4,
  output         io_maskOut_1_1_5,
  output         io_maskOut_1_1_6,
  output         io_maskOut_1_1_7,
  output         io_maskOut_1_1_8,
  output         io_maskOut_1_1_9,
  output         io_maskOut_1_1_10,
  output         io_maskOut_1_1_11,
  output         io_maskOut_1_1_12,
  output         io_maskOut_1_1_13,
  output         io_maskOut_1_1_14,
  output         io_maskOut_1_1_15,
  output         io_maskOut_1_2_0,
  output         io_maskOut_1_2_1,
  output         io_maskOut_1_2_2,
  output         io_maskOut_1_2_3,
  output         io_maskOut_1_2_4,
  output         io_maskOut_1_2_5,
  output         io_maskOut_1_2_6,
  output         io_maskOut_1_2_7,
  output         io_maskOut_1_2_8,
  output         io_maskOut_1_2_9,
  output         io_maskOut_1_2_10,
  output         io_maskOut_1_2_11,
  output         io_maskOut_1_2_12,
  output         io_maskOut_1_2_13,
  output         io_maskOut_1_2_14,
  output         io_maskOut_1_2_15,
  output         io_maskOut_1_3_0,
  output         io_maskOut_1_3_1,
  output         io_maskOut_1_3_2,
  output         io_maskOut_1_3_3,
  output         io_maskOut_1_3_4,
  output         io_maskOut_1_3_5,
  output         io_maskOut_1_3_6,
  output         io_maskOut_1_3_7,
  output         io_maskOut_1_3_8,
  output         io_maskOut_1_3_9,
  output         io_maskOut_1_3_10,
  output         io_maskOut_1_3_11,
  output         io_maskOut_1_3_12,
  output         io_maskOut_1_3_13,
  output         io_maskOut_1_3_14,
  output         io_maskOut_1_3_15,
  output         io_maskOut_2_0_0,
  output         io_maskOut_2_0_1,
  output         io_maskOut_2_0_2,
  output         io_maskOut_2_0_3,
  output         io_maskOut_2_0_4,
  output         io_maskOut_2_0_5,
  output         io_maskOut_2_0_6,
  output         io_maskOut_2_0_7,
  output         io_maskOut_2_0_8,
  output         io_maskOut_2_0_9,
  output         io_maskOut_2_0_10,
  output         io_maskOut_2_0_11,
  output         io_maskOut_2_0_12,
  output         io_maskOut_2_0_13,
  output         io_maskOut_2_0_14,
  output         io_maskOut_2_0_15,
  output         io_maskOut_2_1_0,
  output         io_maskOut_2_1_1,
  output         io_maskOut_2_1_2,
  output         io_maskOut_2_1_3,
  output         io_maskOut_2_1_4,
  output         io_maskOut_2_1_5,
  output         io_maskOut_2_1_6,
  output         io_maskOut_2_1_7,
  output         io_maskOut_2_1_8,
  output         io_maskOut_2_1_9,
  output         io_maskOut_2_1_10,
  output         io_maskOut_2_1_11,
  output         io_maskOut_2_1_12,
  output         io_maskOut_2_1_13,
  output         io_maskOut_2_1_14,
  output         io_maskOut_2_1_15,
  output         io_maskOut_2_2_0,
  output         io_maskOut_2_2_1,
  output         io_maskOut_2_2_2,
  output         io_maskOut_2_2_3,
  output         io_maskOut_2_2_4,
  output         io_maskOut_2_2_5,
  output         io_maskOut_2_2_6,
  output         io_maskOut_2_2_7,
  output         io_maskOut_2_2_8,
  output         io_maskOut_2_2_9,
  output         io_maskOut_2_2_10,
  output         io_maskOut_2_2_11,
  output         io_maskOut_2_2_12,
  output         io_maskOut_2_2_13,
  output         io_maskOut_2_2_14,
  output         io_maskOut_2_2_15,
  output         io_maskOut_2_3_0,
  output         io_maskOut_2_3_1,
  output         io_maskOut_2_3_2,
  output         io_maskOut_2_3_3,
  output         io_maskOut_2_3_4,
  output         io_maskOut_2_3_5,
  output         io_maskOut_2_3_6,
  output         io_maskOut_2_3_7,
  output         io_maskOut_2_3_8,
  output         io_maskOut_2_3_9,
  output         io_maskOut_2_3_10,
  output         io_maskOut_2_3_11,
  output         io_maskOut_2_3_12,
  output         io_maskOut_2_3_13,
  output         io_maskOut_2_3_14,
  output         io_maskOut_2_3_15,
  output         io_maskOut_3_0_0,
  output         io_maskOut_3_0_1,
  output         io_maskOut_3_0_2,
  output         io_maskOut_3_0_3,
  output         io_maskOut_3_0_4,
  output         io_maskOut_3_0_5,
  output         io_maskOut_3_0_6,
  output         io_maskOut_3_0_7,
  output         io_maskOut_3_0_8,
  output         io_maskOut_3_0_9,
  output         io_maskOut_3_0_10,
  output         io_maskOut_3_0_11,
  output         io_maskOut_3_0_12,
  output         io_maskOut_3_0_13,
  output         io_maskOut_3_0_14,
  output         io_maskOut_3_0_15,
  output         io_maskOut_3_1_0,
  output         io_maskOut_3_1_1,
  output         io_maskOut_3_1_2,
  output         io_maskOut_3_1_3,
  output         io_maskOut_3_1_4,
  output         io_maskOut_3_1_5,
  output         io_maskOut_3_1_6,
  output         io_maskOut_3_1_7,
  output         io_maskOut_3_1_8,
  output         io_maskOut_3_1_9,
  output         io_maskOut_3_1_10,
  output         io_maskOut_3_1_11,
  output         io_maskOut_3_1_12,
  output         io_maskOut_3_1_13,
  output         io_maskOut_3_1_14,
  output         io_maskOut_3_1_15,
  output         io_maskOut_3_2_0,
  output         io_maskOut_3_2_1,
  output         io_maskOut_3_2_2,
  output         io_maskOut_3_2_3,
  output         io_maskOut_3_2_4,
  output         io_maskOut_3_2_5,
  output         io_maskOut_3_2_6,
  output         io_maskOut_3_2_7,
  output         io_maskOut_3_2_8,
  output         io_maskOut_3_2_9,
  output         io_maskOut_3_2_10,
  output         io_maskOut_3_2_11,
  output         io_maskOut_3_2_12,
  output         io_maskOut_3_2_13,
  output         io_maskOut_3_2_14,
  output         io_maskOut_3_2_15,
  output         io_maskOut_3_3_0,
  output         io_maskOut_3_3_1,
  output         io_maskOut_3_3_2,
  output         io_maskOut_3_3_3,
  output         io_maskOut_3_3_4,
  output         io_maskOut_3_3_5,
  output         io_maskOut_3_3_6,
  output         io_maskOut_3_3_7,
  output         io_maskOut_3_3_8,
  output         io_maskOut_3_3_9,
  output         io_maskOut_3_3_10,
  output         io_maskOut_3_3_11,
  output         io_maskOut_3_3_12,
  output         io_maskOut_3_3_13,
  output         io_maskOut_3_3_14,
  output         io_maskOut_3_3_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [127:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [127:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [127:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [127:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [127:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [127:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [127:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [127:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] data_0_0_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_0_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_1_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_2_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_0_3_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_0_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_1_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_2_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_1_3_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_0_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_1_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_2_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_2_3_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_0_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_1_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_2_15; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_0; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_1; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_2; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_3; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_4; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_5; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_6; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_7; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_8; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_9; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_10; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_11; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_12; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_13; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_14; // @[Sbuffer.scala 102:17]
  reg [7:0] data_3_3_15; // @[Sbuffer.scala 102:17]
  reg  mask_0_0_0; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_1; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_2; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_3; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_4; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_5; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_6; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_7; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_8; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_9; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_10; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_11; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_12; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_13; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_14; // @[Sbuffer.scala 104:21]
  reg  mask_0_0_15; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_0; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_1; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_2; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_3; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_4; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_5; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_6; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_7; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_8; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_9; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_10; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_11; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_12; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_13; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_14; // @[Sbuffer.scala 104:21]
  reg  mask_0_1_15; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_0; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_1; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_2; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_3; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_4; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_5; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_6; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_7; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_8; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_9; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_10; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_11; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_12; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_13; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_14; // @[Sbuffer.scala 104:21]
  reg  mask_0_2_15; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_0; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_1; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_2; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_3; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_4; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_5; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_6; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_7; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_8; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_9; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_10; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_11; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_12; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_13; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_14; // @[Sbuffer.scala 104:21]
  reg  mask_0_3_15; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_0; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_1; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_2; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_3; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_4; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_5; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_6; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_7; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_8; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_9; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_10; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_11; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_12; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_13; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_14; // @[Sbuffer.scala 104:21]
  reg  mask_1_0_15; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_0; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_1; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_2; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_3; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_4; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_5; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_6; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_7; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_8; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_9; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_10; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_11; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_12; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_13; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_14; // @[Sbuffer.scala 104:21]
  reg  mask_1_1_15; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_0; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_1; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_2; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_3; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_4; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_5; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_6; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_7; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_8; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_9; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_10; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_11; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_12; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_13; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_14; // @[Sbuffer.scala 104:21]
  reg  mask_1_2_15; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_0; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_1; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_2; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_3; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_4; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_5; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_6; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_7; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_8; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_9; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_10; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_11; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_12; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_13; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_14; // @[Sbuffer.scala 104:21]
  reg  mask_1_3_15; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_0; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_1; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_2; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_3; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_4; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_5; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_6; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_7; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_8; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_9; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_10; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_11; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_12; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_13; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_14; // @[Sbuffer.scala 104:21]
  reg  mask_2_0_15; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_0; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_1; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_2; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_3; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_4; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_5; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_6; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_7; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_8; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_9; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_10; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_11; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_12; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_13; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_14; // @[Sbuffer.scala 104:21]
  reg  mask_2_1_15; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_0; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_1; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_2; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_3; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_4; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_5; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_6; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_7; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_8; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_9; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_10; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_11; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_12; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_13; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_14; // @[Sbuffer.scala 104:21]
  reg  mask_2_2_15; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_0; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_1; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_2; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_3; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_4; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_5; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_6; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_7; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_8; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_9; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_10; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_11; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_12; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_13; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_14; // @[Sbuffer.scala 104:21]
  reg  mask_2_3_15; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_0; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_1; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_2; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_3; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_4; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_5; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_6; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_7; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_8; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_9; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_10; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_11; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_12; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_13; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_14; // @[Sbuffer.scala 104:21]
  reg  mask_3_0_15; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_0; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_1; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_2; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_3; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_4; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_5; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_6; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_7; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_8; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_9; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_10; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_11; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_12; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_13; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_14; // @[Sbuffer.scala 104:21]
  reg  mask_3_1_15; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_0; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_1; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_2; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_3; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_4; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_5; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_6; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_7; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_8; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_9; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_10; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_11; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_12; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_13; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_14; // @[Sbuffer.scala 104:21]
  reg  mask_3_2_15; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_0; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_1; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_2; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_3; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_4; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_5; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_6; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_7; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_8; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_9; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_10; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_11; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_12; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_13; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_14; // @[Sbuffer.scala 104:21]
  reg  mask_3_3_15; // @[Sbuffer.scala 104:21]
  reg  line_mask_clean_flag_0; // @[Sbuffer.scala 114:39]
  wire  _GEN_0 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_1 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_2 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_3 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_4 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_5 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_6 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_7 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_8 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_9 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_10 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_11 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_12 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_13 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_14 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_15 = line_mask_clean_flag_0 ? 1'h0 : mask_0_0_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_16 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_17 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_18 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_19 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_20 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_21 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_22 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_23 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_24 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_25 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_26 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_27 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_28 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_29 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_30 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_31 = line_mask_clean_flag_0 ? 1'h0 : mask_0_1_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_32 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_33 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_34 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_35 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_36 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_37 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_38 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_39 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_40 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_41 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_42 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_43 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_44 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_45 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_46 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_47 = line_mask_clean_flag_0 ? 1'h0 : mask_0_2_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_48 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_49 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_50 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_51 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_52 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_53 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_54 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_55 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_56 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_57 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_58 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_59 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_60 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_61 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_62 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_63 = line_mask_clean_flag_0 ? 1'h0 : mask_0_3_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  reg  line_mask_clean_flag_1; // @[Sbuffer.scala 114:39]
  wire  _GEN_64 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_65 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_66 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_67 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_68 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_69 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_70 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_71 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_72 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_73 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_74 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_75 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_76 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_77 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_78 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_79 = line_mask_clean_flag_1 ? 1'h0 : mask_1_0_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_80 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_81 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_82 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_83 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_84 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_85 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_86 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_87 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_88 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_89 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_90 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_91 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_92 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_93 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_94 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_95 = line_mask_clean_flag_1 ? 1'h0 : mask_1_1_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_96 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_97 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_98 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_99 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_100 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_101 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_102 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_103 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_104 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_105 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_106 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_107 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_108 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_109 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_110 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_111 = line_mask_clean_flag_1 ? 1'h0 : mask_1_2_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_112 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_113 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_114 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_115 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_116 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_117 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_118 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_119 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_120 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_121 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_122 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_123 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_124 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_125 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_126 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_127 = line_mask_clean_flag_1 ? 1'h0 : mask_1_3_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  reg  line_mask_clean_flag_2; // @[Sbuffer.scala 114:39]
  wire  _GEN_128 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_129 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_130 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_131 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_132 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_133 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_134 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_135 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_136 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_137 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_138 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_139 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_140 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_141 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_142 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_143 = line_mask_clean_flag_2 ? 1'h0 : mask_2_0_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_144 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_145 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_146 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_147 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_148 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_149 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_150 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_151 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_152 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_153 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_154 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_155 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_156 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_157 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_158 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_159 = line_mask_clean_flag_2 ? 1'h0 : mask_2_1_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_160 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_161 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_162 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_163 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_164 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_165 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_166 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_167 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_168 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_169 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_170 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_171 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_172 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_173 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_174 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_175 = line_mask_clean_flag_2 ? 1'h0 : mask_2_2_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_176 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_177 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_178 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_179 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_180 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_181 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_182 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_183 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_184 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_185 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_186 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_187 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_188 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_189 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_190 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_191 = line_mask_clean_flag_2 ? 1'h0 : mask_2_3_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  reg  line_mask_clean_flag_3; // @[Sbuffer.scala 114:39]
  wire  _GEN_192 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_193 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_194 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_195 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_196 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_197 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_198 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_199 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_200 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_201 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_202 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_203 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_204 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_205 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_206 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_207 = line_mask_clean_flag_3 ? 1'h0 : mask_3_0_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_208 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_209 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_210 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_211 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_212 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_213 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_214 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_215 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_216 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_217 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_218 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_219 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_220 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_221 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_222 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_223 = line_mask_clean_flag_3 ? 1'h0 : mask_3_1_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_224 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_225 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_226 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_227 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_228 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_229 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_230 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_231 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_232 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_233 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_234 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_235 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_236 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_237 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_238 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_239 = line_mask_clean_flag_3 ? 1'h0 : mask_3_2_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_240 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_0; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_241 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_1; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_242 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_2; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_243 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_3; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_244 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_4; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_245 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_5; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_246 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_6; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_247 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_7; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_248 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_8; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_249 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_9; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_250 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_10; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_251 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_11; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_252 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_12; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_253 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_13; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_254 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_14; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  _GEN_255 = line_mask_clean_flag_3 ? 1'h0 : mask_3_3_15; // @[Sbuffer.scala 104:21 118:31 121:34]
  wire  sbuffer_in_s1_line_wen_0 = io_writeReq_0_valid & io_writeReq_0_bits_wvec[0]; // @[Sbuffer.scala 131:46]
  reg  sbuffer_in_s2_line_wen_0; // @[Sbuffer.scala 132:43]
  reg [127:0] line_write_buffer_data_0; // @[Reg.scala 16:16]
  reg  line_write_buffer_wline_0; // @[Reg.scala 16:16]
  reg [15:0] line_write_buffer_mask_0; // @[Reg.scala 16:16]
  reg [1:0] line_write_buffer_offset_0; // @[Reg.scala 16:16]
  wire  _write_byte_T_3 = line_write_buffer_mask_0[0] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte = sbuffer_in_s2_line_wen_0 & _write_byte_T_3; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_7 = line_write_buffer_mask_0[1] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_1 = sbuffer_in_s2_line_wen_0 & _write_byte_T_7; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_11 = line_write_buffer_mask_0[2] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_2 = sbuffer_in_s2_line_wen_0 & _write_byte_T_11; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_15 = line_write_buffer_mask_0[3] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_3 = sbuffer_in_s2_line_wen_0 & _write_byte_T_15; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_19 = line_write_buffer_mask_0[4] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_4 = sbuffer_in_s2_line_wen_0 & _write_byte_T_19; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_23 = line_write_buffer_mask_0[5] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_5 = sbuffer_in_s2_line_wen_0 & _write_byte_T_23; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_27 = line_write_buffer_mask_0[6] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_6 = sbuffer_in_s2_line_wen_0 & _write_byte_T_27; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_31 = line_write_buffer_mask_0[7] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_7 = sbuffer_in_s2_line_wen_0 & _write_byte_T_31; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_35 = line_write_buffer_mask_0[8] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_8 = sbuffer_in_s2_line_wen_0 & _write_byte_T_35; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_39 = line_write_buffer_mask_0[9] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_9 = sbuffer_in_s2_line_wen_0 & _write_byte_T_39; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_43 = line_write_buffer_mask_0[10] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_10 = sbuffer_in_s2_line_wen_0 & _write_byte_T_43; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_47 = line_write_buffer_mask_0[11] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_11 = sbuffer_in_s2_line_wen_0 & _write_byte_T_47; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_51 = line_write_buffer_mask_0[12] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_12 = sbuffer_in_s2_line_wen_0 & _write_byte_T_51; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_55 = line_write_buffer_mask_0[13] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_13 = sbuffer_in_s2_line_wen_0 & _write_byte_T_55; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_59 = line_write_buffer_mask_0[14] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_14 = sbuffer_in_s2_line_wen_0 & _write_byte_T_59; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_63 = line_write_buffer_mask_0[15] & line_write_buffer_offset_0 == 2'h0 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_15 = sbuffer_in_s2_line_wen_0 & _write_byte_T_63; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_67 = line_write_buffer_mask_0[0] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_16 = sbuffer_in_s2_line_wen_0 & _write_byte_T_67; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_71 = line_write_buffer_mask_0[1] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_17 = sbuffer_in_s2_line_wen_0 & _write_byte_T_71; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_75 = line_write_buffer_mask_0[2] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_18 = sbuffer_in_s2_line_wen_0 & _write_byte_T_75; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_79 = line_write_buffer_mask_0[3] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_19 = sbuffer_in_s2_line_wen_0 & _write_byte_T_79; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_83 = line_write_buffer_mask_0[4] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_20 = sbuffer_in_s2_line_wen_0 & _write_byte_T_83; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_87 = line_write_buffer_mask_0[5] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_21 = sbuffer_in_s2_line_wen_0 & _write_byte_T_87; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_91 = line_write_buffer_mask_0[6] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_22 = sbuffer_in_s2_line_wen_0 & _write_byte_T_91; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_95 = line_write_buffer_mask_0[7] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_23 = sbuffer_in_s2_line_wen_0 & _write_byte_T_95; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_99 = line_write_buffer_mask_0[8] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_24 = sbuffer_in_s2_line_wen_0 & _write_byte_T_99; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_103 = line_write_buffer_mask_0[9] & line_write_buffer_offset_0 == 2'h1 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_25 = sbuffer_in_s2_line_wen_0 & _write_byte_T_103; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_107 = line_write_buffer_mask_0[10] & line_write_buffer_offset_0 == 2'h1 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_26 = sbuffer_in_s2_line_wen_0 & _write_byte_T_107; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_111 = line_write_buffer_mask_0[11] & line_write_buffer_offset_0 == 2'h1 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_27 = sbuffer_in_s2_line_wen_0 & _write_byte_T_111; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_115 = line_write_buffer_mask_0[12] & line_write_buffer_offset_0 == 2'h1 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_28 = sbuffer_in_s2_line_wen_0 & _write_byte_T_115; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_119 = line_write_buffer_mask_0[13] & line_write_buffer_offset_0 == 2'h1 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_29 = sbuffer_in_s2_line_wen_0 & _write_byte_T_119; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_123 = line_write_buffer_mask_0[14] & line_write_buffer_offset_0 == 2'h1 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_30 = sbuffer_in_s2_line_wen_0 & _write_byte_T_123; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_127 = line_write_buffer_mask_0[15] & line_write_buffer_offset_0 == 2'h1 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_31 = sbuffer_in_s2_line_wen_0 & _write_byte_T_127; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_131 = line_write_buffer_mask_0[0] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_32 = sbuffer_in_s2_line_wen_0 & _write_byte_T_131; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_135 = line_write_buffer_mask_0[1] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_33 = sbuffer_in_s2_line_wen_0 & _write_byte_T_135; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_139 = line_write_buffer_mask_0[2] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_34 = sbuffer_in_s2_line_wen_0 & _write_byte_T_139; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_143 = line_write_buffer_mask_0[3] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_35 = sbuffer_in_s2_line_wen_0 & _write_byte_T_143; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_147 = line_write_buffer_mask_0[4] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_36 = sbuffer_in_s2_line_wen_0 & _write_byte_T_147; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_151 = line_write_buffer_mask_0[5] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_37 = sbuffer_in_s2_line_wen_0 & _write_byte_T_151; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_155 = line_write_buffer_mask_0[6] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_38 = sbuffer_in_s2_line_wen_0 & _write_byte_T_155; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_159 = line_write_buffer_mask_0[7] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_39 = sbuffer_in_s2_line_wen_0 & _write_byte_T_159; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_163 = line_write_buffer_mask_0[8] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_40 = sbuffer_in_s2_line_wen_0 & _write_byte_T_163; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_167 = line_write_buffer_mask_0[9] & line_write_buffer_offset_0 == 2'h2 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_41 = sbuffer_in_s2_line_wen_0 & _write_byte_T_167; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_171 = line_write_buffer_mask_0[10] & line_write_buffer_offset_0 == 2'h2 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_42 = sbuffer_in_s2_line_wen_0 & _write_byte_T_171; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_175 = line_write_buffer_mask_0[11] & line_write_buffer_offset_0 == 2'h2 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_43 = sbuffer_in_s2_line_wen_0 & _write_byte_T_175; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_179 = line_write_buffer_mask_0[12] & line_write_buffer_offset_0 == 2'h2 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_44 = sbuffer_in_s2_line_wen_0 & _write_byte_T_179; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_183 = line_write_buffer_mask_0[13] & line_write_buffer_offset_0 == 2'h2 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_45 = sbuffer_in_s2_line_wen_0 & _write_byte_T_183; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_187 = line_write_buffer_mask_0[14] & line_write_buffer_offset_0 == 2'h2 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_46 = sbuffer_in_s2_line_wen_0 & _write_byte_T_187; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_191 = line_write_buffer_mask_0[15] & line_write_buffer_offset_0 == 2'h2 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_47 = sbuffer_in_s2_line_wen_0 & _write_byte_T_191; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_195 = line_write_buffer_mask_0[0] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_48 = sbuffer_in_s2_line_wen_0 & _write_byte_T_195; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_199 = line_write_buffer_mask_0[1] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_49 = sbuffer_in_s2_line_wen_0 & _write_byte_T_199; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_203 = line_write_buffer_mask_0[2] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_50 = sbuffer_in_s2_line_wen_0 & _write_byte_T_203; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_207 = line_write_buffer_mask_0[3] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_51 = sbuffer_in_s2_line_wen_0 & _write_byte_T_207; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_211 = line_write_buffer_mask_0[4] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_52 = sbuffer_in_s2_line_wen_0 & _write_byte_T_211; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_215 = line_write_buffer_mask_0[5] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_53 = sbuffer_in_s2_line_wen_0 & _write_byte_T_215; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_219 = line_write_buffer_mask_0[6] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_54 = sbuffer_in_s2_line_wen_0 & _write_byte_T_219; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_223 = line_write_buffer_mask_0[7] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_55 = sbuffer_in_s2_line_wen_0 & _write_byte_T_223; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_227 = line_write_buffer_mask_0[8] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_56 = sbuffer_in_s2_line_wen_0 & _write_byte_T_227; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_231 = line_write_buffer_mask_0[9] & line_write_buffer_offset_0 == 2'h3 | line_write_buffer_wline_0
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_57 = sbuffer_in_s2_line_wen_0 & _write_byte_T_231; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_235 = line_write_buffer_mask_0[10] & line_write_buffer_offset_0 == 2'h3 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_58 = sbuffer_in_s2_line_wen_0 & _write_byte_T_235; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_239 = line_write_buffer_mask_0[11] & line_write_buffer_offset_0 == 2'h3 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_59 = sbuffer_in_s2_line_wen_0 & _write_byte_T_239; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_243 = line_write_buffer_mask_0[12] & line_write_buffer_offset_0 == 2'h3 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_60 = sbuffer_in_s2_line_wen_0 & _write_byte_T_243; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_247 = line_write_buffer_mask_0[13] & line_write_buffer_offset_0 == 2'h3 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_61 = sbuffer_in_s2_line_wen_0 & _write_byte_T_247; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_251 = line_write_buffer_mask_0[14] & line_write_buffer_offset_0 == 2'h3 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_62 = sbuffer_in_s2_line_wen_0 & _write_byte_T_251; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_255 = line_write_buffer_mask_0[15] & line_write_buffer_offset_0 == 2'h3 |
    line_write_buffer_wline_0; // @[Sbuffer.scala 146:83]
  wire  write_byte_63 = sbuffer_in_s2_line_wen_0 & _write_byte_T_255; // @[Sbuffer.scala 145:51]
  wire  sbuffer_in_s1_line_wen_1 = io_writeReq_0_valid & io_writeReq_0_bits_wvec[1]; // @[Sbuffer.scala 131:46]
  reg  sbuffer_in_s2_line_wen_1; // @[Sbuffer.scala 132:43]
  reg [127:0] line_write_buffer_data_1; // @[Reg.scala 16:16]
  reg  line_write_buffer_wline_1; // @[Reg.scala 16:16]
  reg [15:0] line_write_buffer_mask_1; // @[Reg.scala 16:16]
  reg [1:0] line_write_buffer_offset_1; // @[Reg.scala 16:16]
  wire  _write_byte_T_259 = line_write_buffer_mask_1[0] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_64 = sbuffer_in_s2_line_wen_1 & _write_byte_T_259; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_263 = line_write_buffer_mask_1[1] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_65 = sbuffer_in_s2_line_wen_1 & _write_byte_T_263; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_267 = line_write_buffer_mask_1[2] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_66 = sbuffer_in_s2_line_wen_1 & _write_byte_T_267; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_271 = line_write_buffer_mask_1[3] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_67 = sbuffer_in_s2_line_wen_1 & _write_byte_T_271; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_275 = line_write_buffer_mask_1[4] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_68 = sbuffer_in_s2_line_wen_1 & _write_byte_T_275; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_279 = line_write_buffer_mask_1[5] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_69 = sbuffer_in_s2_line_wen_1 & _write_byte_T_279; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_283 = line_write_buffer_mask_1[6] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_70 = sbuffer_in_s2_line_wen_1 & _write_byte_T_283; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_287 = line_write_buffer_mask_1[7] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_71 = sbuffer_in_s2_line_wen_1 & _write_byte_T_287; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_291 = line_write_buffer_mask_1[8] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_72 = sbuffer_in_s2_line_wen_1 & _write_byte_T_291; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_295 = line_write_buffer_mask_1[9] & line_write_buffer_offset_1 == 2'h0 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_73 = sbuffer_in_s2_line_wen_1 & _write_byte_T_295; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_299 = line_write_buffer_mask_1[10] & line_write_buffer_offset_1 == 2'h0 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_74 = sbuffer_in_s2_line_wen_1 & _write_byte_T_299; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_303 = line_write_buffer_mask_1[11] & line_write_buffer_offset_1 == 2'h0 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_75 = sbuffer_in_s2_line_wen_1 & _write_byte_T_303; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_307 = line_write_buffer_mask_1[12] & line_write_buffer_offset_1 == 2'h0 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_76 = sbuffer_in_s2_line_wen_1 & _write_byte_T_307; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_311 = line_write_buffer_mask_1[13] & line_write_buffer_offset_1 == 2'h0 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_77 = sbuffer_in_s2_line_wen_1 & _write_byte_T_311; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_315 = line_write_buffer_mask_1[14] & line_write_buffer_offset_1 == 2'h0 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_78 = sbuffer_in_s2_line_wen_1 & _write_byte_T_315; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_319 = line_write_buffer_mask_1[15] & line_write_buffer_offset_1 == 2'h0 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_79 = sbuffer_in_s2_line_wen_1 & _write_byte_T_319; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_323 = line_write_buffer_mask_1[0] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_80 = sbuffer_in_s2_line_wen_1 & _write_byte_T_323; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_327 = line_write_buffer_mask_1[1] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_81 = sbuffer_in_s2_line_wen_1 & _write_byte_T_327; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_331 = line_write_buffer_mask_1[2] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_82 = sbuffer_in_s2_line_wen_1 & _write_byte_T_331; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_335 = line_write_buffer_mask_1[3] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_83 = sbuffer_in_s2_line_wen_1 & _write_byte_T_335; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_339 = line_write_buffer_mask_1[4] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_84 = sbuffer_in_s2_line_wen_1 & _write_byte_T_339; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_343 = line_write_buffer_mask_1[5] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_85 = sbuffer_in_s2_line_wen_1 & _write_byte_T_343; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_347 = line_write_buffer_mask_1[6] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_86 = sbuffer_in_s2_line_wen_1 & _write_byte_T_347; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_351 = line_write_buffer_mask_1[7] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_87 = sbuffer_in_s2_line_wen_1 & _write_byte_T_351; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_355 = line_write_buffer_mask_1[8] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_88 = sbuffer_in_s2_line_wen_1 & _write_byte_T_355; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_359 = line_write_buffer_mask_1[9] & line_write_buffer_offset_1 == 2'h1 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_89 = sbuffer_in_s2_line_wen_1 & _write_byte_T_359; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_363 = line_write_buffer_mask_1[10] & line_write_buffer_offset_1 == 2'h1 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_90 = sbuffer_in_s2_line_wen_1 & _write_byte_T_363; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_367 = line_write_buffer_mask_1[11] & line_write_buffer_offset_1 == 2'h1 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_91 = sbuffer_in_s2_line_wen_1 & _write_byte_T_367; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_371 = line_write_buffer_mask_1[12] & line_write_buffer_offset_1 == 2'h1 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_92 = sbuffer_in_s2_line_wen_1 & _write_byte_T_371; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_375 = line_write_buffer_mask_1[13] & line_write_buffer_offset_1 == 2'h1 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_93 = sbuffer_in_s2_line_wen_1 & _write_byte_T_375; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_379 = line_write_buffer_mask_1[14] & line_write_buffer_offset_1 == 2'h1 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_94 = sbuffer_in_s2_line_wen_1 & _write_byte_T_379; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_383 = line_write_buffer_mask_1[15] & line_write_buffer_offset_1 == 2'h1 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_95 = sbuffer_in_s2_line_wen_1 & _write_byte_T_383; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_387 = line_write_buffer_mask_1[0] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_96 = sbuffer_in_s2_line_wen_1 & _write_byte_T_387; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_391 = line_write_buffer_mask_1[1] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_97 = sbuffer_in_s2_line_wen_1 & _write_byte_T_391; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_395 = line_write_buffer_mask_1[2] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_98 = sbuffer_in_s2_line_wen_1 & _write_byte_T_395; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_399 = line_write_buffer_mask_1[3] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_99 = sbuffer_in_s2_line_wen_1 & _write_byte_T_399; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_403 = line_write_buffer_mask_1[4] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_100 = sbuffer_in_s2_line_wen_1 & _write_byte_T_403; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_407 = line_write_buffer_mask_1[5] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_101 = sbuffer_in_s2_line_wen_1 & _write_byte_T_407; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_411 = line_write_buffer_mask_1[6] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_102 = sbuffer_in_s2_line_wen_1 & _write_byte_T_411; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_415 = line_write_buffer_mask_1[7] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_103 = sbuffer_in_s2_line_wen_1 & _write_byte_T_415; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_419 = line_write_buffer_mask_1[8] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_104 = sbuffer_in_s2_line_wen_1 & _write_byte_T_419; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_423 = line_write_buffer_mask_1[9] & line_write_buffer_offset_1 == 2'h2 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_105 = sbuffer_in_s2_line_wen_1 & _write_byte_T_423; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_427 = line_write_buffer_mask_1[10] & line_write_buffer_offset_1 == 2'h2 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_106 = sbuffer_in_s2_line_wen_1 & _write_byte_T_427; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_431 = line_write_buffer_mask_1[11] & line_write_buffer_offset_1 == 2'h2 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_107 = sbuffer_in_s2_line_wen_1 & _write_byte_T_431; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_435 = line_write_buffer_mask_1[12] & line_write_buffer_offset_1 == 2'h2 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_108 = sbuffer_in_s2_line_wen_1 & _write_byte_T_435; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_439 = line_write_buffer_mask_1[13] & line_write_buffer_offset_1 == 2'h2 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_109 = sbuffer_in_s2_line_wen_1 & _write_byte_T_439; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_443 = line_write_buffer_mask_1[14] & line_write_buffer_offset_1 == 2'h2 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_110 = sbuffer_in_s2_line_wen_1 & _write_byte_T_443; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_447 = line_write_buffer_mask_1[15] & line_write_buffer_offset_1 == 2'h2 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_111 = sbuffer_in_s2_line_wen_1 & _write_byte_T_447; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_451 = line_write_buffer_mask_1[0] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_112 = sbuffer_in_s2_line_wen_1 & _write_byte_T_451; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_455 = line_write_buffer_mask_1[1] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_113 = sbuffer_in_s2_line_wen_1 & _write_byte_T_455; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_459 = line_write_buffer_mask_1[2] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_114 = sbuffer_in_s2_line_wen_1 & _write_byte_T_459; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_463 = line_write_buffer_mask_1[3] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_115 = sbuffer_in_s2_line_wen_1 & _write_byte_T_463; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_467 = line_write_buffer_mask_1[4] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_116 = sbuffer_in_s2_line_wen_1 & _write_byte_T_467; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_471 = line_write_buffer_mask_1[5] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_117 = sbuffer_in_s2_line_wen_1 & _write_byte_T_471; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_475 = line_write_buffer_mask_1[6] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_118 = sbuffer_in_s2_line_wen_1 & _write_byte_T_475; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_479 = line_write_buffer_mask_1[7] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_119 = sbuffer_in_s2_line_wen_1 & _write_byte_T_479; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_483 = line_write_buffer_mask_1[8] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_120 = sbuffer_in_s2_line_wen_1 & _write_byte_T_483; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_487 = line_write_buffer_mask_1[9] & line_write_buffer_offset_1 == 2'h3 | line_write_buffer_wline_1
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_121 = sbuffer_in_s2_line_wen_1 & _write_byte_T_487; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_491 = line_write_buffer_mask_1[10] & line_write_buffer_offset_1 == 2'h3 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_122 = sbuffer_in_s2_line_wen_1 & _write_byte_T_491; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_495 = line_write_buffer_mask_1[11] & line_write_buffer_offset_1 == 2'h3 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_123 = sbuffer_in_s2_line_wen_1 & _write_byte_T_495; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_499 = line_write_buffer_mask_1[12] & line_write_buffer_offset_1 == 2'h3 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_124 = sbuffer_in_s2_line_wen_1 & _write_byte_T_499; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_503 = line_write_buffer_mask_1[13] & line_write_buffer_offset_1 == 2'h3 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_125 = sbuffer_in_s2_line_wen_1 & _write_byte_T_503; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_507 = line_write_buffer_mask_1[14] & line_write_buffer_offset_1 == 2'h3 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_126 = sbuffer_in_s2_line_wen_1 & _write_byte_T_507; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_511 = line_write_buffer_mask_1[15] & line_write_buffer_offset_1 == 2'h3 |
    line_write_buffer_wline_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_127 = sbuffer_in_s2_line_wen_1 & _write_byte_T_511; // @[Sbuffer.scala 145:51]
  wire  sbuffer_in_s1_line_wen_2 = io_writeReq_0_valid & io_writeReq_0_bits_wvec[2]; // @[Sbuffer.scala 131:46]
  reg  sbuffer_in_s2_line_wen_2; // @[Sbuffer.scala 132:43]
  reg [127:0] line_write_buffer_data_2; // @[Reg.scala 16:16]
  reg  line_write_buffer_wline_2; // @[Reg.scala 16:16]
  reg [15:0] line_write_buffer_mask_2; // @[Reg.scala 16:16]
  reg [1:0] line_write_buffer_offset_2; // @[Reg.scala 16:16]
  wire  _write_byte_T_515 = line_write_buffer_mask_2[0] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_128 = sbuffer_in_s2_line_wen_2 & _write_byte_T_515; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_519 = line_write_buffer_mask_2[1] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_129 = sbuffer_in_s2_line_wen_2 & _write_byte_T_519; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_523 = line_write_buffer_mask_2[2] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_130 = sbuffer_in_s2_line_wen_2 & _write_byte_T_523; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_527 = line_write_buffer_mask_2[3] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_131 = sbuffer_in_s2_line_wen_2 & _write_byte_T_527; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_531 = line_write_buffer_mask_2[4] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_132 = sbuffer_in_s2_line_wen_2 & _write_byte_T_531; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_535 = line_write_buffer_mask_2[5] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_133 = sbuffer_in_s2_line_wen_2 & _write_byte_T_535; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_539 = line_write_buffer_mask_2[6] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_134 = sbuffer_in_s2_line_wen_2 & _write_byte_T_539; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_543 = line_write_buffer_mask_2[7] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_135 = sbuffer_in_s2_line_wen_2 & _write_byte_T_543; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_547 = line_write_buffer_mask_2[8] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_136 = sbuffer_in_s2_line_wen_2 & _write_byte_T_547; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_551 = line_write_buffer_mask_2[9] & line_write_buffer_offset_2 == 2'h0 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_137 = sbuffer_in_s2_line_wen_2 & _write_byte_T_551; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_555 = line_write_buffer_mask_2[10] & line_write_buffer_offset_2 == 2'h0 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_138 = sbuffer_in_s2_line_wen_2 & _write_byte_T_555; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_559 = line_write_buffer_mask_2[11] & line_write_buffer_offset_2 == 2'h0 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_139 = sbuffer_in_s2_line_wen_2 & _write_byte_T_559; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_563 = line_write_buffer_mask_2[12] & line_write_buffer_offset_2 == 2'h0 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_140 = sbuffer_in_s2_line_wen_2 & _write_byte_T_563; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_567 = line_write_buffer_mask_2[13] & line_write_buffer_offset_2 == 2'h0 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_141 = sbuffer_in_s2_line_wen_2 & _write_byte_T_567; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_571 = line_write_buffer_mask_2[14] & line_write_buffer_offset_2 == 2'h0 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_142 = sbuffer_in_s2_line_wen_2 & _write_byte_T_571; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_575 = line_write_buffer_mask_2[15] & line_write_buffer_offset_2 == 2'h0 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_143 = sbuffer_in_s2_line_wen_2 & _write_byte_T_575; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_579 = line_write_buffer_mask_2[0] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_144 = sbuffer_in_s2_line_wen_2 & _write_byte_T_579; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_583 = line_write_buffer_mask_2[1] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_145 = sbuffer_in_s2_line_wen_2 & _write_byte_T_583; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_587 = line_write_buffer_mask_2[2] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_146 = sbuffer_in_s2_line_wen_2 & _write_byte_T_587; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_591 = line_write_buffer_mask_2[3] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_147 = sbuffer_in_s2_line_wen_2 & _write_byte_T_591; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_595 = line_write_buffer_mask_2[4] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_148 = sbuffer_in_s2_line_wen_2 & _write_byte_T_595; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_599 = line_write_buffer_mask_2[5] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_149 = sbuffer_in_s2_line_wen_2 & _write_byte_T_599; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_603 = line_write_buffer_mask_2[6] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_150 = sbuffer_in_s2_line_wen_2 & _write_byte_T_603; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_607 = line_write_buffer_mask_2[7] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_151 = sbuffer_in_s2_line_wen_2 & _write_byte_T_607; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_611 = line_write_buffer_mask_2[8] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_152 = sbuffer_in_s2_line_wen_2 & _write_byte_T_611; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_615 = line_write_buffer_mask_2[9] & line_write_buffer_offset_2 == 2'h1 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_153 = sbuffer_in_s2_line_wen_2 & _write_byte_T_615; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_619 = line_write_buffer_mask_2[10] & line_write_buffer_offset_2 == 2'h1 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_154 = sbuffer_in_s2_line_wen_2 & _write_byte_T_619; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_623 = line_write_buffer_mask_2[11] & line_write_buffer_offset_2 == 2'h1 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_155 = sbuffer_in_s2_line_wen_2 & _write_byte_T_623; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_627 = line_write_buffer_mask_2[12] & line_write_buffer_offset_2 == 2'h1 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_156 = sbuffer_in_s2_line_wen_2 & _write_byte_T_627; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_631 = line_write_buffer_mask_2[13] & line_write_buffer_offset_2 == 2'h1 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_157 = sbuffer_in_s2_line_wen_2 & _write_byte_T_631; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_635 = line_write_buffer_mask_2[14] & line_write_buffer_offset_2 == 2'h1 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_158 = sbuffer_in_s2_line_wen_2 & _write_byte_T_635; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_639 = line_write_buffer_mask_2[15] & line_write_buffer_offset_2 == 2'h1 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_159 = sbuffer_in_s2_line_wen_2 & _write_byte_T_639; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_643 = line_write_buffer_mask_2[0] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_160 = sbuffer_in_s2_line_wen_2 & _write_byte_T_643; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_647 = line_write_buffer_mask_2[1] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_161 = sbuffer_in_s2_line_wen_2 & _write_byte_T_647; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_651 = line_write_buffer_mask_2[2] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_162 = sbuffer_in_s2_line_wen_2 & _write_byte_T_651; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_655 = line_write_buffer_mask_2[3] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_163 = sbuffer_in_s2_line_wen_2 & _write_byte_T_655; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_659 = line_write_buffer_mask_2[4] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_164 = sbuffer_in_s2_line_wen_2 & _write_byte_T_659; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_663 = line_write_buffer_mask_2[5] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_165 = sbuffer_in_s2_line_wen_2 & _write_byte_T_663; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_667 = line_write_buffer_mask_2[6] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_166 = sbuffer_in_s2_line_wen_2 & _write_byte_T_667; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_671 = line_write_buffer_mask_2[7] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_167 = sbuffer_in_s2_line_wen_2 & _write_byte_T_671; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_675 = line_write_buffer_mask_2[8] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_168 = sbuffer_in_s2_line_wen_2 & _write_byte_T_675; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_679 = line_write_buffer_mask_2[9] & line_write_buffer_offset_2 == 2'h2 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_169 = sbuffer_in_s2_line_wen_2 & _write_byte_T_679; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_683 = line_write_buffer_mask_2[10] & line_write_buffer_offset_2 == 2'h2 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_170 = sbuffer_in_s2_line_wen_2 & _write_byte_T_683; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_687 = line_write_buffer_mask_2[11] & line_write_buffer_offset_2 == 2'h2 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_171 = sbuffer_in_s2_line_wen_2 & _write_byte_T_687; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_691 = line_write_buffer_mask_2[12] & line_write_buffer_offset_2 == 2'h2 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_172 = sbuffer_in_s2_line_wen_2 & _write_byte_T_691; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_695 = line_write_buffer_mask_2[13] & line_write_buffer_offset_2 == 2'h2 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_173 = sbuffer_in_s2_line_wen_2 & _write_byte_T_695; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_699 = line_write_buffer_mask_2[14] & line_write_buffer_offset_2 == 2'h2 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_174 = sbuffer_in_s2_line_wen_2 & _write_byte_T_699; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_703 = line_write_buffer_mask_2[15] & line_write_buffer_offset_2 == 2'h2 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_175 = sbuffer_in_s2_line_wen_2 & _write_byte_T_703; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_707 = line_write_buffer_mask_2[0] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_176 = sbuffer_in_s2_line_wen_2 & _write_byte_T_707; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_711 = line_write_buffer_mask_2[1] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_177 = sbuffer_in_s2_line_wen_2 & _write_byte_T_711; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_715 = line_write_buffer_mask_2[2] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_178 = sbuffer_in_s2_line_wen_2 & _write_byte_T_715; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_719 = line_write_buffer_mask_2[3] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_179 = sbuffer_in_s2_line_wen_2 & _write_byte_T_719; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_723 = line_write_buffer_mask_2[4] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_180 = sbuffer_in_s2_line_wen_2 & _write_byte_T_723; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_727 = line_write_buffer_mask_2[5] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_181 = sbuffer_in_s2_line_wen_2 & _write_byte_T_727; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_731 = line_write_buffer_mask_2[6] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_182 = sbuffer_in_s2_line_wen_2 & _write_byte_T_731; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_735 = line_write_buffer_mask_2[7] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_183 = sbuffer_in_s2_line_wen_2 & _write_byte_T_735; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_739 = line_write_buffer_mask_2[8] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_184 = sbuffer_in_s2_line_wen_2 & _write_byte_T_739; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_743 = line_write_buffer_mask_2[9] & line_write_buffer_offset_2 == 2'h3 | line_write_buffer_wline_2
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_185 = sbuffer_in_s2_line_wen_2 & _write_byte_T_743; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_747 = line_write_buffer_mask_2[10] & line_write_buffer_offset_2 == 2'h3 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_186 = sbuffer_in_s2_line_wen_2 & _write_byte_T_747; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_751 = line_write_buffer_mask_2[11] & line_write_buffer_offset_2 == 2'h3 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_187 = sbuffer_in_s2_line_wen_2 & _write_byte_T_751; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_755 = line_write_buffer_mask_2[12] & line_write_buffer_offset_2 == 2'h3 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_188 = sbuffer_in_s2_line_wen_2 & _write_byte_T_755; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_759 = line_write_buffer_mask_2[13] & line_write_buffer_offset_2 == 2'h3 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_189 = sbuffer_in_s2_line_wen_2 & _write_byte_T_759; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_763 = line_write_buffer_mask_2[14] & line_write_buffer_offset_2 == 2'h3 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_190 = sbuffer_in_s2_line_wen_2 & _write_byte_T_763; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_767 = line_write_buffer_mask_2[15] & line_write_buffer_offset_2 == 2'h3 |
    line_write_buffer_wline_2; // @[Sbuffer.scala 146:83]
  wire  write_byte_191 = sbuffer_in_s2_line_wen_2 & _write_byte_T_767; // @[Sbuffer.scala 145:51]
  wire  sbuffer_in_s1_line_wen_3 = io_writeReq_0_valid & io_writeReq_0_bits_wvec[3]; // @[Sbuffer.scala 131:46]
  reg  sbuffer_in_s2_line_wen_3; // @[Sbuffer.scala 132:43]
  reg [127:0] line_write_buffer_data_3; // @[Reg.scala 16:16]
  reg  line_write_buffer_wline_3; // @[Reg.scala 16:16]
  reg [15:0] line_write_buffer_mask_3; // @[Reg.scala 16:16]
  reg [1:0] line_write_buffer_offset_3; // @[Reg.scala 16:16]
  wire  _write_byte_T_771 = line_write_buffer_mask_3[0] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_192 = sbuffer_in_s2_line_wen_3 & _write_byte_T_771; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_775 = line_write_buffer_mask_3[1] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_193 = sbuffer_in_s2_line_wen_3 & _write_byte_T_775; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_779 = line_write_buffer_mask_3[2] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_194 = sbuffer_in_s2_line_wen_3 & _write_byte_T_779; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_783 = line_write_buffer_mask_3[3] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_195 = sbuffer_in_s2_line_wen_3 & _write_byte_T_783; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_787 = line_write_buffer_mask_3[4] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_196 = sbuffer_in_s2_line_wen_3 & _write_byte_T_787; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_791 = line_write_buffer_mask_3[5] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_197 = sbuffer_in_s2_line_wen_3 & _write_byte_T_791; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_795 = line_write_buffer_mask_3[6] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_198 = sbuffer_in_s2_line_wen_3 & _write_byte_T_795; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_799 = line_write_buffer_mask_3[7] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_199 = sbuffer_in_s2_line_wen_3 & _write_byte_T_799; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_803 = line_write_buffer_mask_3[8] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_200 = sbuffer_in_s2_line_wen_3 & _write_byte_T_803; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_807 = line_write_buffer_mask_3[9] & line_write_buffer_offset_3 == 2'h0 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_201 = sbuffer_in_s2_line_wen_3 & _write_byte_T_807; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_811 = line_write_buffer_mask_3[10] & line_write_buffer_offset_3 == 2'h0 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_202 = sbuffer_in_s2_line_wen_3 & _write_byte_T_811; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_815 = line_write_buffer_mask_3[11] & line_write_buffer_offset_3 == 2'h0 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_203 = sbuffer_in_s2_line_wen_3 & _write_byte_T_815; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_819 = line_write_buffer_mask_3[12] & line_write_buffer_offset_3 == 2'h0 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_204 = sbuffer_in_s2_line_wen_3 & _write_byte_T_819; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_823 = line_write_buffer_mask_3[13] & line_write_buffer_offset_3 == 2'h0 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_205 = sbuffer_in_s2_line_wen_3 & _write_byte_T_823; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_827 = line_write_buffer_mask_3[14] & line_write_buffer_offset_3 == 2'h0 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_206 = sbuffer_in_s2_line_wen_3 & _write_byte_T_827; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_831 = line_write_buffer_mask_3[15] & line_write_buffer_offset_3 == 2'h0 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_207 = sbuffer_in_s2_line_wen_3 & _write_byte_T_831; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_835 = line_write_buffer_mask_3[0] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_208 = sbuffer_in_s2_line_wen_3 & _write_byte_T_835; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_839 = line_write_buffer_mask_3[1] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_209 = sbuffer_in_s2_line_wen_3 & _write_byte_T_839; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_843 = line_write_buffer_mask_3[2] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_210 = sbuffer_in_s2_line_wen_3 & _write_byte_T_843; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_847 = line_write_buffer_mask_3[3] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_211 = sbuffer_in_s2_line_wen_3 & _write_byte_T_847; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_851 = line_write_buffer_mask_3[4] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_212 = sbuffer_in_s2_line_wen_3 & _write_byte_T_851; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_855 = line_write_buffer_mask_3[5] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_213 = sbuffer_in_s2_line_wen_3 & _write_byte_T_855; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_859 = line_write_buffer_mask_3[6] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_214 = sbuffer_in_s2_line_wen_3 & _write_byte_T_859; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_863 = line_write_buffer_mask_3[7] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_215 = sbuffer_in_s2_line_wen_3 & _write_byte_T_863; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_867 = line_write_buffer_mask_3[8] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_216 = sbuffer_in_s2_line_wen_3 & _write_byte_T_867; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_871 = line_write_buffer_mask_3[9] & line_write_buffer_offset_3 == 2'h1 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_217 = sbuffer_in_s2_line_wen_3 & _write_byte_T_871; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_875 = line_write_buffer_mask_3[10] & line_write_buffer_offset_3 == 2'h1 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_218 = sbuffer_in_s2_line_wen_3 & _write_byte_T_875; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_879 = line_write_buffer_mask_3[11] & line_write_buffer_offset_3 == 2'h1 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_219 = sbuffer_in_s2_line_wen_3 & _write_byte_T_879; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_883 = line_write_buffer_mask_3[12] & line_write_buffer_offset_3 == 2'h1 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_220 = sbuffer_in_s2_line_wen_3 & _write_byte_T_883; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_887 = line_write_buffer_mask_3[13] & line_write_buffer_offset_3 == 2'h1 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_221 = sbuffer_in_s2_line_wen_3 & _write_byte_T_887; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_891 = line_write_buffer_mask_3[14] & line_write_buffer_offset_3 == 2'h1 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_222 = sbuffer_in_s2_line_wen_3 & _write_byte_T_891; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_895 = line_write_buffer_mask_3[15] & line_write_buffer_offset_3 == 2'h1 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_223 = sbuffer_in_s2_line_wen_3 & _write_byte_T_895; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_899 = line_write_buffer_mask_3[0] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_224 = sbuffer_in_s2_line_wen_3 & _write_byte_T_899; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_903 = line_write_buffer_mask_3[1] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_225 = sbuffer_in_s2_line_wen_3 & _write_byte_T_903; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_907 = line_write_buffer_mask_3[2] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_226 = sbuffer_in_s2_line_wen_3 & _write_byte_T_907; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_911 = line_write_buffer_mask_3[3] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_227 = sbuffer_in_s2_line_wen_3 & _write_byte_T_911; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_915 = line_write_buffer_mask_3[4] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_228 = sbuffer_in_s2_line_wen_3 & _write_byte_T_915; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_919 = line_write_buffer_mask_3[5] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_229 = sbuffer_in_s2_line_wen_3 & _write_byte_T_919; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_923 = line_write_buffer_mask_3[6] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_230 = sbuffer_in_s2_line_wen_3 & _write_byte_T_923; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_927 = line_write_buffer_mask_3[7] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_231 = sbuffer_in_s2_line_wen_3 & _write_byte_T_927; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_931 = line_write_buffer_mask_3[8] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_232 = sbuffer_in_s2_line_wen_3 & _write_byte_T_931; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_935 = line_write_buffer_mask_3[9] & line_write_buffer_offset_3 == 2'h2 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_233 = sbuffer_in_s2_line_wen_3 & _write_byte_T_935; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_939 = line_write_buffer_mask_3[10] & line_write_buffer_offset_3 == 2'h2 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_234 = sbuffer_in_s2_line_wen_3 & _write_byte_T_939; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_943 = line_write_buffer_mask_3[11] & line_write_buffer_offset_3 == 2'h2 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_235 = sbuffer_in_s2_line_wen_3 & _write_byte_T_943; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_947 = line_write_buffer_mask_3[12] & line_write_buffer_offset_3 == 2'h2 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_236 = sbuffer_in_s2_line_wen_3 & _write_byte_T_947; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_951 = line_write_buffer_mask_3[13] & line_write_buffer_offset_3 == 2'h2 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_237 = sbuffer_in_s2_line_wen_3 & _write_byte_T_951; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_955 = line_write_buffer_mask_3[14] & line_write_buffer_offset_3 == 2'h2 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_238 = sbuffer_in_s2_line_wen_3 & _write_byte_T_955; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_959 = line_write_buffer_mask_3[15] & line_write_buffer_offset_3 == 2'h2 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_239 = sbuffer_in_s2_line_wen_3 & _write_byte_T_959; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_963 = line_write_buffer_mask_3[0] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_240 = sbuffer_in_s2_line_wen_3 & _write_byte_T_963; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_967 = line_write_buffer_mask_3[1] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_241 = sbuffer_in_s2_line_wen_3 & _write_byte_T_967; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_971 = line_write_buffer_mask_3[2] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_242 = sbuffer_in_s2_line_wen_3 & _write_byte_T_971; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_975 = line_write_buffer_mask_3[3] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_243 = sbuffer_in_s2_line_wen_3 & _write_byte_T_975; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_979 = line_write_buffer_mask_3[4] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_244 = sbuffer_in_s2_line_wen_3 & _write_byte_T_979; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_983 = line_write_buffer_mask_3[5] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_245 = sbuffer_in_s2_line_wen_3 & _write_byte_T_983; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_987 = line_write_buffer_mask_3[6] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_246 = sbuffer_in_s2_line_wen_3 & _write_byte_T_987; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_991 = line_write_buffer_mask_3[7] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_247 = sbuffer_in_s2_line_wen_3 & _write_byte_T_991; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_995 = line_write_buffer_mask_3[8] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_248 = sbuffer_in_s2_line_wen_3 & _write_byte_T_995; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_999 = line_write_buffer_mask_3[9] & line_write_buffer_offset_3 == 2'h3 | line_write_buffer_wline_3
    ; // @[Sbuffer.scala 146:83]
  wire  write_byte_249 = sbuffer_in_s2_line_wen_3 & _write_byte_T_999; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1003 = line_write_buffer_mask_3[10] & line_write_buffer_offset_3 == 2'h3 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_250 = sbuffer_in_s2_line_wen_3 & _write_byte_T_1003; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1007 = line_write_buffer_mask_3[11] & line_write_buffer_offset_3 == 2'h3 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_251 = sbuffer_in_s2_line_wen_3 & _write_byte_T_1007; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1011 = line_write_buffer_mask_3[12] & line_write_buffer_offset_3 == 2'h3 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_252 = sbuffer_in_s2_line_wen_3 & _write_byte_T_1011; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1015 = line_write_buffer_mask_3[13] & line_write_buffer_offset_3 == 2'h3 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_253 = sbuffer_in_s2_line_wen_3 & _write_byte_T_1015; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1019 = line_write_buffer_mask_3[14] & line_write_buffer_offset_3 == 2'h3 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_254 = sbuffer_in_s2_line_wen_3 & _write_byte_T_1019; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1023 = line_write_buffer_mask_3[15] & line_write_buffer_offset_3 == 2'h3 |
    line_write_buffer_wline_3; // @[Sbuffer.scala 146:83]
  wire  write_byte_255 = sbuffer_in_s2_line_wen_3 & _write_byte_T_1023; // @[Sbuffer.scala 145:51]
  wire  sbuffer_in_s1_line_wen_0_1 = io_writeReq_1_valid & io_writeReq_1_bits_wvec[0]; // @[Sbuffer.scala 131:46]
  reg  sbuffer_in_s2_line_wen_0_1; // @[Sbuffer.scala 132:43]
  reg [127:0] line_write_buffer_data_0_1; // @[Reg.scala 16:16]
  reg  line_write_buffer_wline_0_1; // @[Reg.scala 16:16]
  reg [15:0] line_write_buffer_mask_0_1; // @[Reg.scala 16:16]
  reg [1:0] line_write_buffer_offset_0_1; // @[Reg.scala 16:16]
  wire  _write_byte_T_1027 = line_write_buffer_mask_0_1[0] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_256 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1027; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1031 = line_write_buffer_mask_0_1[1] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_257 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1031; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1035 = line_write_buffer_mask_0_1[2] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_258 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1035; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1039 = line_write_buffer_mask_0_1[3] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_259 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1039; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1043 = line_write_buffer_mask_0_1[4] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_260 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1043; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1047 = line_write_buffer_mask_0_1[5] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_261 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1047; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1051 = line_write_buffer_mask_0_1[6] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_262 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1051; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1055 = line_write_buffer_mask_0_1[7] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_263 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1055; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1059 = line_write_buffer_mask_0_1[8] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_264 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1059; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1063 = line_write_buffer_mask_0_1[9] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_265 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1063; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1067 = line_write_buffer_mask_0_1[10] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_266 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1067; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1071 = line_write_buffer_mask_0_1[11] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_267 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1071; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1075 = line_write_buffer_mask_0_1[12] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_268 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1075; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1079 = line_write_buffer_mask_0_1[13] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_269 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1079; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1083 = line_write_buffer_mask_0_1[14] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_270 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1083; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1087 = line_write_buffer_mask_0_1[15] & line_write_buffer_offset_0_1 == 2'h0 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_271 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1087; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1091 = line_write_buffer_mask_0_1[0] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_272 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1091; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1095 = line_write_buffer_mask_0_1[1] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_273 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1095; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1099 = line_write_buffer_mask_0_1[2] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_274 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1099; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1103 = line_write_buffer_mask_0_1[3] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_275 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1103; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1107 = line_write_buffer_mask_0_1[4] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_276 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1107; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1111 = line_write_buffer_mask_0_1[5] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_277 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1111; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1115 = line_write_buffer_mask_0_1[6] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_278 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1115; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1119 = line_write_buffer_mask_0_1[7] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_279 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1119; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1123 = line_write_buffer_mask_0_1[8] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_280 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1123; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1127 = line_write_buffer_mask_0_1[9] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_281 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1127; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1131 = line_write_buffer_mask_0_1[10] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_282 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1131; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1135 = line_write_buffer_mask_0_1[11] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_283 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1135; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1139 = line_write_buffer_mask_0_1[12] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_284 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1139; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1143 = line_write_buffer_mask_0_1[13] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_285 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1143; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1147 = line_write_buffer_mask_0_1[14] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_286 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1147; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1151 = line_write_buffer_mask_0_1[15] & line_write_buffer_offset_0_1 == 2'h1 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_287 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1151; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1155 = line_write_buffer_mask_0_1[0] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_288 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1155; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1159 = line_write_buffer_mask_0_1[1] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_289 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1159; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1163 = line_write_buffer_mask_0_1[2] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_290 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1163; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1167 = line_write_buffer_mask_0_1[3] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_291 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1167; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1171 = line_write_buffer_mask_0_1[4] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_292 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1171; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1175 = line_write_buffer_mask_0_1[5] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_293 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1175; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1179 = line_write_buffer_mask_0_1[6] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_294 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1179; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1183 = line_write_buffer_mask_0_1[7] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_295 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1183; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1187 = line_write_buffer_mask_0_1[8] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_296 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1187; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1191 = line_write_buffer_mask_0_1[9] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_297 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1191; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1195 = line_write_buffer_mask_0_1[10] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_298 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1195; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1199 = line_write_buffer_mask_0_1[11] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_299 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1199; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1203 = line_write_buffer_mask_0_1[12] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_300 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1203; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1207 = line_write_buffer_mask_0_1[13] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_301 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1207; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1211 = line_write_buffer_mask_0_1[14] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_302 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1211; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1215 = line_write_buffer_mask_0_1[15] & line_write_buffer_offset_0_1 == 2'h2 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_303 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1215; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1219 = line_write_buffer_mask_0_1[0] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_304 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1219; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1223 = line_write_buffer_mask_0_1[1] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_305 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1223; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1227 = line_write_buffer_mask_0_1[2] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_306 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1227; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1231 = line_write_buffer_mask_0_1[3] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_307 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1231; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1235 = line_write_buffer_mask_0_1[4] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_308 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1235; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1239 = line_write_buffer_mask_0_1[5] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_309 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1239; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1243 = line_write_buffer_mask_0_1[6] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_310 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1243; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1247 = line_write_buffer_mask_0_1[7] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_311 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1247; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1251 = line_write_buffer_mask_0_1[8] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_312 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1251; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1255 = line_write_buffer_mask_0_1[9] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_313 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1255; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1259 = line_write_buffer_mask_0_1[10] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_314 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1259; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1263 = line_write_buffer_mask_0_1[11] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_315 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1263; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1267 = line_write_buffer_mask_0_1[12] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_316 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1267; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1271 = line_write_buffer_mask_0_1[13] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_317 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1271; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1275 = line_write_buffer_mask_0_1[14] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_318 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1275; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1279 = line_write_buffer_mask_0_1[15] & line_write_buffer_offset_0_1 == 2'h3 |
    line_write_buffer_wline_0_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_319 = sbuffer_in_s2_line_wen_0_1 & _write_byte_T_1279; // @[Sbuffer.scala 145:51]
  wire  sbuffer_in_s1_line_wen_1_1 = io_writeReq_1_valid & io_writeReq_1_bits_wvec[1]; // @[Sbuffer.scala 131:46]
  reg  sbuffer_in_s2_line_wen_1_1; // @[Sbuffer.scala 132:43]
  reg [127:0] line_write_buffer_data_1_1; // @[Reg.scala 16:16]
  reg  line_write_buffer_wline_1_1; // @[Reg.scala 16:16]
  reg [15:0] line_write_buffer_mask_1_1; // @[Reg.scala 16:16]
  reg [1:0] line_write_buffer_offset_1_1; // @[Reg.scala 16:16]
  wire  _write_byte_T_1283 = line_write_buffer_mask_1_1[0] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_320 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1283; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1287 = line_write_buffer_mask_1_1[1] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_321 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1287; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1291 = line_write_buffer_mask_1_1[2] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_322 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1291; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1295 = line_write_buffer_mask_1_1[3] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_323 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1295; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1299 = line_write_buffer_mask_1_1[4] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_324 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1299; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1303 = line_write_buffer_mask_1_1[5] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_325 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1303; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1307 = line_write_buffer_mask_1_1[6] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_326 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1307; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1311 = line_write_buffer_mask_1_1[7] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_327 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1311; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1315 = line_write_buffer_mask_1_1[8] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_328 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1315; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1319 = line_write_buffer_mask_1_1[9] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_329 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1319; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1323 = line_write_buffer_mask_1_1[10] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_330 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1323; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1327 = line_write_buffer_mask_1_1[11] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_331 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1327; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1331 = line_write_buffer_mask_1_1[12] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_332 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1331; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1335 = line_write_buffer_mask_1_1[13] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_333 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1335; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1339 = line_write_buffer_mask_1_1[14] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_334 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1339; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1343 = line_write_buffer_mask_1_1[15] & line_write_buffer_offset_1_1 == 2'h0 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_335 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1343; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1347 = line_write_buffer_mask_1_1[0] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_336 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1347; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1351 = line_write_buffer_mask_1_1[1] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_337 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1351; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1355 = line_write_buffer_mask_1_1[2] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_338 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1355; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1359 = line_write_buffer_mask_1_1[3] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_339 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1359; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1363 = line_write_buffer_mask_1_1[4] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_340 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1363; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1367 = line_write_buffer_mask_1_1[5] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_341 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1367; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1371 = line_write_buffer_mask_1_1[6] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_342 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1371; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1375 = line_write_buffer_mask_1_1[7] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_343 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1375; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1379 = line_write_buffer_mask_1_1[8] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_344 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1379; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1383 = line_write_buffer_mask_1_1[9] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_345 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1383; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1387 = line_write_buffer_mask_1_1[10] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_346 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1387; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1391 = line_write_buffer_mask_1_1[11] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_347 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1391; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1395 = line_write_buffer_mask_1_1[12] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_348 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1395; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1399 = line_write_buffer_mask_1_1[13] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_349 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1399; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1403 = line_write_buffer_mask_1_1[14] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_350 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1403; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1407 = line_write_buffer_mask_1_1[15] & line_write_buffer_offset_1_1 == 2'h1 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_351 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1407; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1411 = line_write_buffer_mask_1_1[0] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_352 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1411; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1415 = line_write_buffer_mask_1_1[1] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_353 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1415; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1419 = line_write_buffer_mask_1_1[2] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_354 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1419; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1423 = line_write_buffer_mask_1_1[3] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_355 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1423; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1427 = line_write_buffer_mask_1_1[4] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_356 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1427; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1431 = line_write_buffer_mask_1_1[5] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_357 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1431; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1435 = line_write_buffer_mask_1_1[6] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_358 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1435; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1439 = line_write_buffer_mask_1_1[7] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_359 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1439; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1443 = line_write_buffer_mask_1_1[8] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_360 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1443; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1447 = line_write_buffer_mask_1_1[9] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_361 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1447; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1451 = line_write_buffer_mask_1_1[10] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_362 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1451; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1455 = line_write_buffer_mask_1_1[11] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_363 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1455; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1459 = line_write_buffer_mask_1_1[12] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_364 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1459; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1463 = line_write_buffer_mask_1_1[13] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_365 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1463; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1467 = line_write_buffer_mask_1_1[14] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_366 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1467; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1471 = line_write_buffer_mask_1_1[15] & line_write_buffer_offset_1_1 == 2'h2 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_367 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1471; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1475 = line_write_buffer_mask_1_1[0] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_368 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1475; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1479 = line_write_buffer_mask_1_1[1] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_369 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1479; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1483 = line_write_buffer_mask_1_1[2] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_370 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1483; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1487 = line_write_buffer_mask_1_1[3] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_371 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1487; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1491 = line_write_buffer_mask_1_1[4] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_372 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1491; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1495 = line_write_buffer_mask_1_1[5] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_373 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1495; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1499 = line_write_buffer_mask_1_1[6] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_374 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1499; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1503 = line_write_buffer_mask_1_1[7] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_375 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1503; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1507 = line_write_buffer_mask_1_1[8] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_376 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1507; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1511 = line_write_buffer_mask_1_1[9] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_377 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1511; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1515 = line_write_buffer_mask_1_1[10] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_378 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1515; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1519 = line_write_buffer_mask_1_1[11] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_379 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1519; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1523 = line_write_buffer_mask_1_1[12] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_380 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1523; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1527 = line_write_buffer_mask_1_1[13] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_381 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1527; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1531 = line_write_buffer_mask_1_1[14] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_382 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1531; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1535 = line_write_buffer_mask_1_1[15] & line_write_buffer_offset_1_1 == 2'h3 |
    line_write_buffer_wline_1_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_383 = sbuffer_in_s2_line_wen_1_1 & _write_byte_T_1535; // @[Sbuffer.scala 145:51]
  wire  sbuffer_in_s1_line_wen_2_1 = io_writeReq_1_valid & io_writeReq_1_bits_wvec[2]; // @[Sbuffer.scala 131:46]
  reg  sbuffer_in_s2_line_wen_2_1; // @[Sbuffer.scala 132:43]
  reg [127:0] line_write_buffer_data_2_1; // @[Reg.scala 16:16]
  reg  line_write_buffer_wline_2_1; // @[Reg.scala 16:16]
  reg [15:0] line_write_buffer_mask_2_1; // @[Reg.scala 16:16]
  reg [1:0] line_write_buffer_offset_2_1; // @[Reg.scala 16:16]
  wire  _write_byte_T_1539 = line_write_buffer_mask_2_1[0] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_384 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1539; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1543 = line_write_buffer_mask_2_1[1] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_385 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1543; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1547 = line_write_buffer_mask_2_1[2] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_386 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1547; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1551 = line_write_buffer_mask_2_1[3] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_387 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1551; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1555 = line_write_buffer_mask_2_1[4] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_388 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1555; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1559 = line_write_buffer_mask_2_1[5] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_389 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1559; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1563 = line_write_buffer_mask_2_1[6] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_390 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1563; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1567 = line_write_buffer_mask_2_1[7] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_391 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1567; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1571 = line_write_buffer_mask_2_1[8] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_392 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1571; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1575 = line_write_buffer_mask_2_1[9] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_393 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1575; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1579 = line_write_buffer_mask_2_1[10] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_394 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1579; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1583 = line_write_buffer_mask_2_1[11] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_395 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1583; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1587 = line_write_buffer_mask_2_1[12] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_396 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1587; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1591 = line_write_buffer_mask_2_1[13] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_397 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1591; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1595 = line_write_buffer_mask_2_1[14] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_398 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1595; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1599 = line_write_buffer_mask_2_1[15] & line_write_buffer_offset_2_1 == 2'h0 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_399 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1599; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1603 = line_write_buffer_mask_2_1[0] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_400 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1603; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1607 = line_write_buffer_mask_2_1[1] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_401 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1607; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1611 = line_write_buffer_mask_2_1[2] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_402 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1611; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1615 = line_write_buffer_mask_2_1[3] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_403 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1615; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1619 = line_write_buffer_mask_2_1[4] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_404 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1619; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1623 = line_write_buffer_mask_2_1[5] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_405 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1623; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1627 = line_write_buffer_mask_2_1[6] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_406 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1627; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1631 = line_write_buffer_mask_2_1[7] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_407 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1631; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1635 = line_write_buffer_mask_2_1[8] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_408 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1635; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1639 = line_write_buffer_mask_2_1[9] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_409 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1639; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1643 = line_write_buffer_mask_2_1[10] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_410 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1643; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1647 = line_write_buffer_mask_2_1[11] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_411 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1647; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1651 = line_write_buffer_mask_2_1[12] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_412 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1651; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1655 = line_write_buffer_mask_2_1[13] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_413 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1655; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1659 = line_write_buffer_mask_2_1[14] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_414 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1659; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1663 = line_write_buffer_mask_2_1[15] & line_write_buffer_offset_2_1 == 2'h1 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_415 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1663; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1667 = line_write_buffer_mask_2_1[0] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_416 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1667; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1671 = line_write_buffer_mask_2_1[1] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_417 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1671; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1675 = line_write_buffer_mask_2_1[2] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_418 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1675; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1679 = line_write_buffer_mask_2_1[3] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_419 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1679; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1683 = line_write_buffer_mask_2_1[4] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_420 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1683; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1687 = line_write_buffer_mask_2_1[5] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_421 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1687; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1691 = line_write_buffer_mask_2_1[6] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_422 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1691; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1695 = line_write_buffer_mask_2_1[7] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_423 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1695; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1699 = line_write_buffer_mask_2_1[8] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_424 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1699; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1703 = line_write_buffer_mask_2_1[9] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_425 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1703; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1707 = line_write_buffer_mask_2_1[10] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_426 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1707; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1711 = line_write_buffer_mask_2_1[11] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_427 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1711; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1715 = line_write_buffer_mask_2_1[12] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_428 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1715; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1719 = line_write_buffer_mask_2_1[13] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_429 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1719; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1723 = line_write_buffer_mask_2_1[14] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_430 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1723; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1727 = line_write_buffer_mask_2_1[15] & line_write_buffer_offset_2_1 == 2'h2 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_431 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1727; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1731 = line_write_buffer_mask_2_1[0] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_432 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1731; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1735 = line_write_buffer_mask_2_1[1] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_433 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1735; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1739 = line_write_buffer_mask_2_1[2] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_434 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1739; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1743 = line_write_buffer_mask_2_1[3] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_435 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1743; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1747 = line_write_buffer_mask_2_1[4] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_436 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1747; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1751 = line_write_buffer_mask_2_1[5] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_437 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1751; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1755 = line_write_buffer_mask_2_1[6] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_438 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1755; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1759 = line_write_buffer_mask_2_1[7] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_439 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1759; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1763 = line_write_buffer_mask_2_1[8] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_440 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1763; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1767 = line_write_buffer_mask_2_1[9] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_441 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1767; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1771 = line_write_buffer_mask_2_1[10] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_442 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1771; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1775 = line_write_buffer_mask_2_1[11] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_443 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1775; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1779 = line_write_buffer_mask_2_1[12] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_444 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1779; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1783 = line_write_buffer_mask_2_1[13] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_445 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1783; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1787 = line_write_buffer_mask_2_1[14] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_446 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1787; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1791 = line_write_buffer_mask_2_1[15] & line_write_buffer_offset_2_1 == 2'h3 |
    line_write_buffer_wline_2_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_447 = sbuffer_in_s2_line_wen_2_1 & _write_byte_T_1791; // @[Sbuffer.scala 145:51]
  wire  sbuffer_in_s1_line_wen_3_1 = io_writeReq_1_valid & io_writeReq_1_bits_wvec[3]; // @[Sbuffer.scala 131:46]
  reg  sbuffer_in_s2_line_wen_3_1; // @[Sbuffer.scala 132:43]
  reg [127:0] line_write_buffer_data_3_1; // @[Reg.scala 16:16]
  reg  line_write_buffer_wline_3_1; // @[Reg.scala 16:16]
  reg [15:0] line_write_buffer_mask_3_1; // @[Reg.scala 16:16]
  reg [1:0] line_write_buffer_offset_3_1; // @[Reg.scala 16:16]
  wire  _write_byte_T_1795 = line_write_buffer_mask_3_1[0] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_448 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1795; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1799 = line_write_buffer_mask_3_1[1] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_449 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1799; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1803 = line_write_buffer_mask_3_1[2] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_450 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1803; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1807 = line_write_buffer_mask_3_1[3] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_451 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1807; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1811 = line_write_buffer_mask_3_1[4] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_452 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1811; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1815 = line_write_buffer_mask_3_1[5] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_453 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1815; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1819 = line_write_buffer_mask_3_1[6] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_454 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1819; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1823 = line_write_buffer_mask_3_1[7] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_455 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1823; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1827 = line_write_buffer_mask_3_1[8] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_456 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1827; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1831 = line_write_buffer_mask_3_1[9] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_457 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1831; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1835 = line_write_buffer_mask_3_1[10] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_458 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1835; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1839 = line_write_buffer_mask_3_1[11] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_459 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1839; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1843 = line_write_buffer_mask_3_1[12] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_460 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1843; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1847 = line_write_buffer_mask_3_1[13] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_461 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1847; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1851 = line_write_buffer_mask_3_1[14] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_462 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1851; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1855 = line_write_buffer_mask_3_1[15] & line_write_buffer_offset_3_1 == 2'h0 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_463 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1855; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1859 = line_write_buffer_mask_3_1[0] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_464 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1859; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1863 = line_write_buffer_mask_3_1[1] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_465 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1863; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1867 = line_write_buffer_mask_3_1[2] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_466 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1867; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1871 = line_write_buffer_mask_3_1[3] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_467 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1871; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1875 = line_write_buffer_mask_3_1[4] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_468 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1875; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1879 = line_write_buffer_mask_3_1[5] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_469 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1879; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1883 = line_write_buffer_mask_3_1[6] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_470 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1883; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1887 = line_write_buffer_mask_3_1[7] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_471 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1887; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1891 = line_write_buffer_mask_3_1[8] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_472 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1891; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1895 = line_write_buffer_mask_3_1[9] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_473 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1895; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1899 = line_write_buffer_mask_3_1[10] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_474 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1899; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1903 = line_write_buffer_mask_3_1[11] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_475 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1903; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1907 = line_write_buffer_mask_3_1[12] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_476 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1907; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1911 = line_write_buffer_mask_3_1[13] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_477 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1911; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1915 = line_write_buffer_mask_3_1[14] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_478 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1915; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1919 = line_write_buffer_mask_3_1[15] & line_write_buffer_offset_3_1 == 2'h1 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_479 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1919; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1923 = line_write_buffer_mask_3_1[0] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_480 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1923; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1927 = line_write_buffer_mask_3_1[1] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_481 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1927; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1931 = line_write_buffer_mask_3_1[2] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_482 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1931; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1935 = line_write_buffer_mask_3_1[3] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_483 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1935; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1939 = line_write_buffer_mask_3_1[4] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_484 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1939; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1943 = line_write_buffer_mask_3_1[5] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_485 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1943; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1947 = line_write_buffer_mask_3_1[6] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_486 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1947; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1951 = line_write_buffer_mask_3_1[7] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_487 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1951; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1955 = line_write_buffer_mask_3_1[8] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_488 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1955; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1959 = line_write_buffer_mask_3_1[9] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_489 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1959; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1963 = line_write_buffer_mask_3_1[10] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_490 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1963; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1967 = line_write_buffer_mask_3_1[11] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_491 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1967; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1971 = line_write_buffer_mask_3_1[12] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_492 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1971; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1975 = line_write_buffer_mask_3_1[13] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_493 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1975; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1979 = line_write_buffer_mask_3_1[14] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_494 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1979; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1983 = line_write_buffer_mask_3_1[15] & line_write_buffer_offset_3_1 == 2'h2 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_495 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1983; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1987 = line_write_buffer_mask_3_1[0] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_496 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1987; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1991 = line_write_buffer_mask_3_1[1] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_497 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1991; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1995 = line_write_buffer_mask_3_1[2] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_498 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1995; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_1999 = line_write_buffer_mask_3_1[3] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_499 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_1999; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2003 = line_write_buffer_mask_3_1[4] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_500 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2003; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2007 = line_write_buffer_mask_3_1[5] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_501 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2007; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2011 = line_write_buffer_mask_3_1[6] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_502 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2011; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2015 = line_write_buffer_mask_3_1[7] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_503 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2015; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2019 = line_write_buffer_mask_3_1[8] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_504 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2019; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2023 = line_write_buffer_mask_3_1[9] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_505 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2023; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2027 = line_write_buffer_mask_3_1[10] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_506 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2027; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2031 = line_write_buffer_mask_3_1[11] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_507 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2031; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2035 = line_write_buffer_mask_3_1[12] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_508 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2035; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2039 = line_write_buffer_mask_3_1[13] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_509 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2039; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2043 = line_write_buffer_mask_3_1[14] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_510 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2043; // @[Sbuffer.scala 145:51]
  wire  _write_byte_T_2047 = line_write_buffer_mask_3_1[15] & line_write_buffer_offset_3_1 == 2'h3 |
    line_write_buffer_wline_3_1; // @[Sbuffer.scala 146:83]
  wire  write_byte_511 = sbuffer_in_s2_line_wen_3_1 & _write_byte_T_2047; // @[Sbuffer.scala 145:51]
  assign io_dataOut_0_0_0 = data_0_0_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_1 = data_0_0_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_2 = data_0_0_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_3 = data_0_0_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_4 = data_0_0_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_5 = data_0_0_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_6 = data_0_0_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_7 = data_0_0_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_8 = data_0_0_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_9 = data_0_0_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_10 = data_0_0_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_11 = data_0_0_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_12 = data_0_0_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_13 = data_0_0_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_14 = data_0_0_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_0_15 = data_0_0_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_0 = data_0_1_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_1 = data_0_1_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_2 = data_0_1_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_3 = data_0_1_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_4 = data_0_1_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_5 = data_0_1_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_6 = data_0_1_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_7 = data_0_1_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_8 = data_0_1_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_9 = data_0_1_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_10 = data_0_1_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_11 = data_0_1_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_12 = data_0_1_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_13 = data_0_1_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_14 = data_0_1_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_1_15 = data_0_1_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_0 = data_0_2_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_1 = data_0_2_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_2 = data_0_2_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_3 = data_0_2_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_4 = data_0_2_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_5 = data_0_2_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_6 = data_0_2_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_7 = data_0_2_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_8 = data_0_2_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_9 = data_0_2_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_10 = data_0_2_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_11 = data_0_2_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_12 = data_0_2_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_13 = data_0_2_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_14 = data_0_2_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_2_15 = data_0_2_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_0 = data_0_3_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_1 = data_0_3_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_2 = data_0_3_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_3 = data_0_3_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_4 = data_0_3_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_5 = data_0_3_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_6 = data_0_3_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_7 = data_0_3_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_8 = data_0_3_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_9 = data_0_3_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_10 = data_0_3_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_11 = data_0_3_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_12 = data_0_3_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_13 = data_0_3_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_14 = data_0_3_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_0_3_15 = data_0_3_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_0 = data_1_0_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_1 = data_1_0_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_2 = data_1_0_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_3 = data_1_0_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_4 = data_1_0_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_5 = data_1_0_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_6 = data_1_0_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_7 = data_1_0_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_8 = data_1_0_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_9 = data_1_0_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_10 = data_1_0_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_11 = data_1_0_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_12 = data_1_0_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_13 = data_1_0_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_14 = data_1_0_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_0_15 = data_1_0_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_0 = data_1_1_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_1 = data_1_1_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_2 = data_1_1_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_3 = data_1_1_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_4 = data_1_1_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_5 = data_1_1_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_6 = data_1_1_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_7 = data_1_1_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_8 = data_1_1_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_9 = data_1_1_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_10 = data_1_1_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_11 = data_1_1_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_12 = data_1_1_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_13 = data_1_1_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_14 = data_1_1_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_1_15 = data_1_1_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_0 = data_1_2_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_1 = data_1_2_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_2 = data_1_2_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_3 = data_1_2_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_4 = data_1_2_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_5 = data_1_2_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_6 = data_1_2_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_7 = data_1_2_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_8 = data_1_2_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_9 = data_1_2_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_10 = data_1_2_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_11 = data_1_2_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_12 = data_1_2_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_13 = data_1_2_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_14 = data_1_2_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_2_15 = data_1_2_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_0 = data_1_3_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_1 = data_1_3_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_2 = data_1_3_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_3 = data_1_3_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_4 = data_1_3_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_5 = data_1_3_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_6 = data_1_3_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_7 = data_1_3_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_8 = data_1_3_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_9 = data_1_3_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_10 = data_1_3_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_11 = data_1_3_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_12 = data_1_3_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_13 = data_1_3_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_14 = data_1_3_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_1_3_15 = data_1_3_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_0 = data_2_0_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_1 = data_2_0_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_2 = data_2_0_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_3 = data_2_0_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_4 = data_2_0_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_5 = data_2_0_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_6 = data_2_0_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_7 = data_2_0_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_8 = data_2_0_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_9 = data_2_0_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_10 = data_2_0_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_11 = data_2_0_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_12 = data_2_0_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_13 = data_2_0_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_14 = data_2_0_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_0_15 = data_2_0_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_0 = data_2_1_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_1 = data_2_1_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_2 = data_2_1_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_3 = data_2_1_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_4 = data_2_1_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_5 = data_2_1_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_6 = data_2_1_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_7 = data_2_1_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_8 = data_2_1_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_9 = data_2_1_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_10 = data_2_1_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_11 = data_2_1_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_12 = data_2_1_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_13 = data_2_1_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_14 = data_2_1_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_1_15 = data_2_1_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_0 = data_2_2_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_1 = data_2_2_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_2 = data_2_2_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_3 = data_2_2_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_4 = data_2_2_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_5 = data_2_2_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_6 = data_2_2_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_7 = data_2_2_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_8 = data_2_2_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_9 = data_2_2_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_10 = data_2_2_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_11 = data_2_2_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_12 = data_2_2_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_13 = data_2_2_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_14 = data_2_2_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_2_15 = data_2_2_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_0 = data_2_3_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_1 = data_2_3_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_2 = data_2_3_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_3 = data_2_3_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_4 = data_2_3_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_5 = data_2_3_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_6 = data_2_3_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_7 = data_2_3_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_8 = data_2_3_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_9 = data_2_3_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_10 = data_2_3_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_11 = data_2_3_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_12 = data_2_3_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_13 = data_2_3_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_14 = data_2_3_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_2_3_15 = data_2_3_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_0 = data_3_0_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_1 = data_3_0_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_2 = data_3_0_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_3 = data_3_0_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_4 = data_3_0_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_5 = data_3_0_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_6 = data_3_0_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_7 = data_3_0_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_8 = data_3_0_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_9 = data_3_0_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_10 = data_3_0_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_11 = data_3_0_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_12 = data_3_0_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_13 = data_3_0_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_14 = data_3_0_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_0_15 = data_3_0_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_0 = data_3_1_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_1 = data_3_1_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_2 = data_3_1_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_3 = data_3_1_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_4 = data_3_1_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_5 = data_3_1_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_6 = data_3_1_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_7 = data_3_1_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_8 = data_3_1_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_9 = data_3_1_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_10 = data_3_1_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_11 = data_3_1_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_12 = data_3_1_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_13 = data_3_1_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_14 = data_3_1_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_1_15 = data_3_1_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_0 = data_3_2_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_1 = data_3_2_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_2 = data_3_2_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_3 = data_3_2_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_4 = data_3_2_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_5 = data_3_2_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_6 = data_3_2_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_7 = data_3_2_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_8 = data_3_2_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_9 = data_3_2_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_10 = data_3_2_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_11 = data_3_2_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_12 = data_3_2_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_13 = data_3_2_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_14 = data_3_2_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_2_15 = data_3_2_15; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_0 = data_3_3_0; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_1 = data_3_3_1; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_2 = data_3_3_2; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_3 = data_3_3_3; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_4 = data_3_3_4; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_5 = data_3_3_5; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_6 = data_3_3_6; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_7 = data_3_3_7; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_8 = data_3_3_8; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_9 = data_3_3_9; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_10 = data_3_3_10; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_11 = data_3_3_11; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_12 = data_3_3_12; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_13 = data_3_3_13; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_14 = data_3_3_14; // @[Sbuffer.scala 182:14]
  assign io_dataOut_3_3_15 = data_3_3_15; // @[Sbuffer.scala 182:14]
  assign io_maskOut_0_0_0 = mask_0_0_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_1 = mask_0_0_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_2 = mask_0_0_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_3 = mask_0_0_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_4 = mask_0_0_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_5 = mask_0_0_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_6 = mask_0_0_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_7 = mask_0_0_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_8 = mask_0_0_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_9 = mask_0_0_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_10 = mask_0_0_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_11 = mask_0_0_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_12 = mask_0_0_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_13 = mask_0_0_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_14 = mask_0_0_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_0_15 = mask_0_0_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_0 = mask_0_1_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_1 = mask_0_1_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_2 = mask_0_1_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_3 = mask_0_1_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_4 = mask_0_1_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_5 = mask_0_1_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_6 = mask_0_1_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_7 = mask_0_1_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_8 = mask_0_1_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_9 = mask_0_1_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_10 = mask_0_1_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_11 = mask_0_1_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_12 = mask_0_1_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_13 = mask_0_1_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_14 = mask_0_1_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_1_15 = mask_0_1_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_0 = mask_0_2_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_1 = mask_0_2_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_2 = mask_0_2_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_3 = mask_0_2_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_4 = mask_0_2_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_5 = mask_0_2_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_6 = mask_0_2_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_7 = mask_0_2_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_8 = mask_0_2_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_9 = mask_0_2_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_10 = mask_0_2_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_11 = mask_0_2_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_12 = mask_0_2_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_13 = mask_0_2_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_14 = mask_0_2_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_2_15 = mask_0_2_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_0 = mask_0_3_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_1 = mask_0_3_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_2 = mask_0_3_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_3 = mask_0_3_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_4 = mask_0_3_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_5 = mask_0_3_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_6 = mask_0_3_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_7 = mask_0_3_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_8 = mask_0_3_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_9 = mask_0_3_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_10 = mask_0_3_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_11 = mask_0_3_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_12 = mask_0_3_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_13 = mask_0_3_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_14 = mask_0_3_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_0_3_15 = mask_0_3_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_0 = mask_1_0_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_1 = mask_1_0_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_2 = mask_1_0_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_3 = mask_1_0_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_4 = mask_1_0_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_5 = mask_1_0_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_6 = mask_1_0_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_7 = mask_1_0_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_8 = mask_1_0_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_9 = mask_1_0_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_10 = mask_1_0_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_11 = mask_1_0_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_12 = mask_1_0_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_13 = mask_1_0_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_14 = mask_1_0_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_0_15 = mask_1_0_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_0 = mask_1_1_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_1 = mask_1_1_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_2 = mask_1_1_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_3 = mask_1_1_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_4 = mask_1_1_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_5 = mask_1_1_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_6 = mask_1_1_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_7 = mask_1_1_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_8 = mask_1_1_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_9 = mask_1_1_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_10 = mask_1_1_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_11 = mask_1_1_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_12 = mask_1_1_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_13 = mask_1_1_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_14 = mask_1_1_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_1_15 = mask_1_1_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_0 = mask_1_2_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_1 = mask_1_2_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_2 = mask_1_2_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_3 = mask_1_2_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_4 = mask_1_2_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_5 = mask_1_2_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_6 = mask_1_2_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_7 = mask_1_2_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_8 = mask_1_2_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_9 = mask_1_2_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_10 = mask_1_2_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_11 = mask_1_2_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_12 = mask_1_2_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_13 = mask_1_2_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_14 = mask_1_2_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_2_15 = mask_1_2_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_0 = mask_1_3_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_1 = mask_1_3_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_2 = mask_1_3_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_3 = mask_1_3_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_4 = mask_1_3_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_5 = mask_1_3_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_6 = mask_1_3_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_7 = mask_1_3_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_8 = mask_1_3_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_9 = mask_1_3_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_10 = mask_1_3_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_11 = mask_1_3_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_12 = mask_1_3_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_13 = mask_1_3_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_14 = mask_1_3_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_1_3_15 = mask_1_3_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_0 = mask_2_0_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_1 = mask_2_0_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_2 = mask_2_0_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_3 = mask_2_0_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_4 = mask_2_0_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_5 = mask_2_0_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_6 = mask_2_0_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_7 = mask_2_0_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_8 = mask_2_0_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_9 = mask_2_0_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_10 = mask_2_0_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_11 = mask_2_0_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_12 = mask_2_0_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_13 = mask_2_0_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_14 = mask_2_0_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_0_15 = mask_2_0_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_0 = mask_2_1_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_1 = mask_2_1_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_2 = mask_2_1_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_3 = mask_2_1_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_4 = mask_2_1_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_5 = mask_2_1_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_6 = mask_2_1_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_7 = mask_2_1_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_8 = mask_2_1_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_9 = mask_2_1_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_10 = mask_2_1_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_11 = mask_2_1_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_12 = mask_2_1_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_13 = mask_2_1_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_14 = mask_2_1_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_1_15 = mask_2_1_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_0 = mask_2_2_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_1 = mask_2_2_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_2 = mask_2_2_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_3 = mask_2_2_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_4 = mask_2_2_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_5 = mask_2_2_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_6 = mask_2_2_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_7 = mask_2_2_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_8 = mask_2_2_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_9 = mask_2_2_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_10 = mask_2_2_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_11 = mask_2_2_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_12 = mask_2_2_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_13 = mask_2_2_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_14 = mask_2_2_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_2_15 = mask_2_2_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_0 = mask_2_3_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_1 = mask_2_3_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_2 = mask_2_3_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_3 = mask_2_3_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_4 = mask_2_3_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_5 = mask_2_3_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_6 = mask_2_3_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_7 = mask_2_3_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_8 = mask_2_3_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_9 = mask_2_3_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_10 = mask_2_3_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_11 = mask_2_3_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_12 = mask_2_3_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_13 = mask_2_3_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_14 = mask_2_3_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_2_3_15 = mask_2_3_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_0 = mask_3_0_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_1 = mask_3_0_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_2 = mask_3_0_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_3 = mask_3_0_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_4 = mask_3_0_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_5 = mask_3_0_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_6 = mask_3_0_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_7 = mask_3_0_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_8 = mask_3_0_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_9 = mask_3_0_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_10 = mask_3_0_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_11 = mask_3_0_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_12 = mask_3_0_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_13 = mask_3_0_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_14 = mask_3_0_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_0_15 = mask_3_0_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_0 = mask_3_1_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_1 = mask_3_1_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_2 = mask_3_1_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_3 = mask_3_1_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_4 = mask_3_1_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_5 = mask_3_1_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_6 = mask_3_1_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_7 = mask_3_1_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_8 = mask_3_1_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_9 = mask_3_1_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_10 = mask_3_1_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_11 = mask_3_1_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_12 = mask_3_1_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_13 = mask_3_1_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_14 = mask_3_1_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_1_15 = mask_3_1_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_0 = mask_3_2_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_1 = mask_3_2_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_2 = mask_3_2_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_3 = mask_3_2_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_4 = mask_3_2_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_5 = mask_3_2_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_6 = mask_3_2_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_7 = mask_3_2_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_8 = mask_3_2_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_9 = mask_3_2_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_10 = mask_3_2_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_11 = mask_3_2_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_12 = mask_3_2_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_13 = mask_3_2_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_14 = mask_3_2_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_2_15 = mask_3_2_15; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_0 = mask_3_3_0; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_1 = mask_3_3_1; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_2 = mask_3_3_2; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_3 = mask_3_3_3; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_4 = mask_3_3_4; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_5 = mask_3_3_5; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_6 = mask_3_3_6; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_7 = mask_3_3_7; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_8 = mask_3_3_8; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_9 = mask_3_3_9; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_10 = mask_3_3_10; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_11 = mask_3_3_11; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_12 = mask_3_3_12; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_13 = mask_3_3_13; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_14 = mask_3_3_14; // @[Sbuffer.scala 183:14]
  assign io_maskOut_3_3_15 = mask_3_3_15; // @[Sbuffer.scala 183:14]
  always @(posedge clock) begin
    if (write_byte_256) begin // @[Sbuffer.scala 149:27]
      data_0_0_0 <= line_write_buffer_data_0_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte) begin // @[Sbuffer.scala 149:27]
      data_0_0_0 <= line_write_buffer_data_0[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_257) begin // @[Sbuffer.scala 149:27]
      data_0_0_1 <= line_write_buffer_data_0_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_1) begin // @[Sbuffer.scala 149:27]
      data_0_0_1 <= line_write_buffer_data_0[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_258) begin // @[Sbuffer.scala 149:27]
      data_0_0_2 <= line_write_buffer_data_0_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_2) begin // @[Sbuffer.scala 149:27]
      data_0_0_2 <= line_write_buffer_data_0[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_259) begin // @[Sbuffer.scala 149:27]
      data_0_0_3 <= line_write_buffer_data_0_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_3) begin // @[Sbuffer.scala 149:27]
      data_0_0_3 <= line_write_buffer_data_0[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_260) begin // @[Sbuffer.scala 149:27]
      data_0_0_4 <= line_write_buffer_data_0_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_4) begin // @[Sbuffer.scala 149:27]
      data_0_0_4 <= line_write_buffer_data_0[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_261) begin // @[Sbuffer.scala 149:27]
      data_0_0_5 <= line_write_buffer_data_0_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_5) begin // @[Sbuffer.scala 149:27]
      data_0_0_5 <= line_write_buffer_data_0[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_262) begin // @[Sbuffer.scala 149:27]
      data_0_0_6 <= line_write_buffer_data_0_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_6) begin // @[Sbuffer.scala 149:27]
      data_0_0_6 <= line_write_buffer_data_0[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_263) begin // @[Sbuffer.scala 149:27]
      data_0_0_7 <= line_write_buffer_data_0_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_7) begin // @[Sbuffer.scala 149:27]
      data_0_0_7 <= line_write_buffer_data_0[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_264) begin // @[Sbuffer.scala 149:27]
      data_0_0_8 <= line_write_buffer_data_0_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_8) begin // @[Sbuffer.scala 149:27]
      data_0_0_8 <= line_write_buffer_data_0[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_265) begin // @[Sbuffer.scala 149:27]
      data_0_0_9 <= line_write_buffer_data_0_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_9) begin // @[Sbuffer.scala 149:27]
      data_0_0_9 <= line_write_buffer_data_0[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_266) begin // @[Sbuffer.scala 149:27]
      data_0_0_10 <= line_write_buffer_data_0_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_10) begin // @[Sbuffer.scala 149:27]
      data_0_0_10 <= line_write_buffer_data_0[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_267) begin // @[Sbuffer.scala 149:27]
      data_0_0_11 <= line_write_buffer_data_0_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_11) begin // @[Sbuffer.scala 149:27]
      data_0_0_11 <= line_write_buffer_data_0[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_268) begin // @[Sbuffer.scala 149:27]
      data_0_0_12 <= line_write_buffer_data_0_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_12) begin // @[Sbuffer.scala 149:27]
      data_0_0_12 <= line_write_buffer_data_0[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_269) begin // @[Sbuffer.scala 149:27]
      data_0_0_13 <= line_write_buffer_data_0_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_13) begin // @[Sbuffer.scala 149:27]
      data_0_0_13 <= line_write_buffer_data_0[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_270) begin // @[Sbuffer.scala 149:27]
      data_0_0_14 <= line_write_buffer_data_0_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_14) begin // @[Sbuffer.scala 149:27]
      data_0_0_14 <= line_write_buffer_data_0[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_271) begin // @[Sbuffer.scala 149:27]
      data_0_0_15 <= line_write_buffer_data_0_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_15) begin // @[Sbuffer.scala 149:27]
      data_0_0_15 <= line_write_buffer_data_0[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_272) begin // @[Sbuffer.scala 149:27]
      data_0_1_0 <= line_write_buffer_data_0_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_16) begin // @[Sbuffer.scala 149:27]
      data_0_1_0 <= line_write_buffer_data_0[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_273) begin // @[Sbuffer.scala 149:27]
      data_0_1_1 <= line_write_buffer_data_0_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_17) begin // @[Sbuffer.scala 149:27]
      data_0_1_1 <= line_write_buffer_data_0[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_274) begin // @[Sbuffer.scala 149:27]
      data_0_1_2 <= line_write_buffer_data_0_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_18) begin // @[Sbuffer.scala 149:27]
      data_0_1_2 <= line_write_buffer_data_0[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_275) begin // @[Sbuffer.scala 149:27]
      data_0_1_3 <= line_write_buffer_data_0_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_19) begin // @[Sbuffer.scala 149:27]
      data_0_1_3 <= line_write_buffer_data_0[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_276) begin // @[Sbuffer.scala 149:27]
      data_0_1_4 <= line_write_buffer_data_0_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_20) begin // @[Sbuffer.scala 149:27]
      data_0_1_4 <= line_write_buffer_data_0[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_277) begin // @[Sbuffer.scala 149:27]
      data_0_1_5 <= line_write_buffer_data_0_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_21) begin // @[Sbuffer.scala 149:27]
      data_0_1_5 <= line_write_buffer_data_0[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_278) begin // @[Sbuffer.scala 149:27]
      data_0_1_6 <= line_write_buffer_data_0_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_22) begin // @[Sbuffer.scala 149:27]
      data_0_1_6 <= line_write_buffer_data_0[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_279) begin // @[Sbuffer.scala 149:27]
      data_0_1_7 <= line_write_buffer_data_0_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_23) begin // @[Sbuffer.scala 149:27]
      data_0_1_7 <= line_write_buffer_data_0[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_280) begin // @[Sbuffer.scala 149:27]
      data_0_1_8 <= line_write_buffer_data_0_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_24) begin // @[Sbuffer.scala 149:27]
      data_0_1_8 <= line_write_buffer_data_0[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_281) begin // @[Sbuffer.scala 149:27]
      data_0_1_9 <= line_write_buffer_data_0_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_25) begin // @[Sbuffer.scala 149:27]
      data_0_1_9 <= line_write_buffer_data_0[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_282) begin // @[Sbuffer.scala 149:27]
      data_0_1_10 <= line_write_buffer_data_0_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_26) begin // @[Sbuffer.scala 149:27]
      data_0_1_10 <= line_write_buffer_data_0[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_283) begin // @[Sbuffer.scala 149:27]
      data_0_1_11 <= line_write_buffer_data_0_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_27) begin // @[Sbuffer.scala 149:27]
      data_0_1_11 <= line_write_buffer_data_0[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_284) begin // @[Sbuffer.scala 149:27]
      data_0_1_12 <= line_write_buffer_data_0_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_28) begin // @[Sbuffer.scala 149:27]
      data_0_1_12 <= line_write_buffer_data_0[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_285) begin // @[Sbuffer.scala 149:27]
      data_0_1_13 <= line_write_buffer_data_0_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_29) begin // @[Sbuffer.scala 149:27]
      data_0_1_13 <= line_write_buffer_data_0[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_286) begin // @[Sbuffer.scala 149:27]
      data_0_1_14 <= line_write_buffer_data_0_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_30) begin // @[Sbuffer.scala 149:27]
      data_0_1_14 <= line_write_buffer_data_0[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_287) begin // @[Sbuffer.scala 149:27]
      data_0_1_15 <= line_write_buffer_data_0_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_31) begin // @[Sbuffer.scala 149:27]
      data_0_1_15 <= line_write_buffer_data_0[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_288) begin // @[Sbuffer.scala 149:27]
      data_0_2_0 <= line_write_buffer_data_0_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_32) begin // @[Sbuffer.scala 149:27]
      data_0_2_0 <= line_write_buffer_data_0[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_289) begin // @[Sbuffer.scala 149:27]
      data_0_2_1 <= line_write_buffer_data_0_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_33) begin // @[Sbuffer.scala 149:27]
      data_0_2_1 <= line_write_buffer_data_0[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_290) begin // @[Sbuffer.scala 149:27]
      data_0_2_2 <= line_write_buffer_data_0_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_34) begin // @[Sbuffer.scala 149:27]
      data_0_2_2 <= line_write_buffer_data_0[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_291) begin // @[Sbuffer.scala 149:27]
      data_0_2_3 <= line_write_buffer_data_0_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_35) begin // @[Sbuffer.scala 149:27]
      data_0_2_3 <= line_write_buffer_data_0[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_292) begin // @[Sbuffer.scala 149:27]
      data_0_2_4 <= line_write_buffer_data_0_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_36) begin // @[Sbuffer.scala 149:27]
      data_0_2_4 <= line_write_buffer_data_0[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_293) begin // @[Sbuffer.scala 149:27]
      data_0_2_5 <= line_write_buffer_data_0_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_37) begin // @[Sbuffer.scala 149:27]
      data_0_2_5 <= line_write_buffer_data_0[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_294) begin // @[Sbuffer.scala 149:27]
      data_0_2_6 <= line_write_buffer_data_0_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_38) begin // @[Sbuffer.scala 149:27]
      data_0_2_6 <= line_write_buffer_data_0[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_295) begin // @[Sbuffer.scala 149:27]
      data_0_2_7 <= line_write_buffer_data_0_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_39) begin // @[Sbuffer.scala 149:27]
      data_0_2_7 <= line_write_buffer_data_0[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_296) begin // @[Sbuffer.scala 149:27]
      data_0_2_8 <= line_write_buffer_data_0_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_40) begin // @[Sbuffer.scala 149:27]
      data_0_2_8 <= line_write_buffer_data_0[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_297) begin // @[Sbuffer.scala 149:27]
      data_0_2_9 <= line_write_buffer_data_0_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_41) begin // @[Sbuffer.scala 149:27]
      data_0_2_9 <= line_write_buffer_data_0[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_298) begin // @[Sbuffer.scala 149:27]
      data_0_2_10 <= line_write_buffer_data_0_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_42) begin // @[Sbuffer.scala 149:27]
      data_0_2_10 <= line_write_buffer_data_0[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_299) begin // @[Sbuffer.scala 149:27]
      data_0_2_11 <= line_write_buffer_data_0_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_43) begin // @[Sbuffer.scala 149:27]
      data_0_2_11 <= line_write_buffer_data_0[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_300) begin // @[Sbuffer.scala 149:27]
      data_0_2_12 <= line_write_buffer_data_0_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_44) begin // @[Sbuffer.scala 149:27]
      data_0_2_12 <= line_write_buffer_data_0[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_301) begin // @[Sbuffer.scala 149:27]
      data_0_2_13 <= line_write_buffer_data_0_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_45) begin // @[Sbuffer.scala 149:27]
      data_0_2_13 <= line_write_buffer_data_0[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_302) begin // @[Sbuffer.scala 149:27]
      data_0_2_14 <= line_write_buffer_data_0_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_46) begin // @[Sbuffer.scala 149:27]
      data_0_2_14 <= line_write_buffer_data_0[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_303) begin // @[Sbuffer.scala 149:27]
      data_0_2_15 <= line_write_buffer_data_0_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_47) begin // @[Sbuffer.scala 149:27]
      data_0_2_15 <= line_write_buffer_data_0[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_304) begin // @[Sbuffer.scala 149:27]
      data_0_3_0 <= line_write_buffer_data_0_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_48) begin // @[Sbuffer.scala 149:27]
      data_0_3_0 <= line_write_buffer_data_0[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_305) begin // @[Sbuffer.scala 149:27]
      data_0_3_1 <= line_write_buffer_data_0_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_49) begin // @[Sbuffer.scala 149:27]
      data_0_3_1 <= line_write_buffer_data_0[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_306) begin // @[Sbuffer.scala 149:27]
      data_0_3_2 <= line_write_buffer_data_0_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_50) begin // @[Sbuffer.scala 149:27]
      data_0_3_2 <= line_write_buffer_data_0[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_307) begin // @[Sbuffer.scala 149:27]
      data_0_3_3 <= line_write_buffer_data_0_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_51) begin // @[Sbuffer.scala 149:27]
      data_0_3_3 <= line_write_buffer_data_0[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_308) begin // @[Sbuffer.scala 149:27]
      data_0_3_4 <= line_write_buffer_data_0_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_52) begin // @[Sbuffer.scala 149:27]
      data_0_3_4 <= line_write_buffer_data_0[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_309) begin // @[Sbuffer.scala 149:27]
      data_0_3_5 <= line_write_buffer_data_0_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_53) begin // @[Sbuffer.scala 149:27]
      data_0_3_5 <= line_write_buffer_data_0[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_310) begin // @[Sbuffer.scala 149:27]
      data_0_3_6 <= line_write_buffer_data_0_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_54) begin // @[Sbuffer.scala 149:27]
      data_0_3_6 <= line_write_buffer_data_0[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_311) begin // @[Sbuffer.scala 149:27]
      data_0_3_7 <= line_write_buffer_data_0_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_55) begin // @[Sbuffer.scala 149:27]
      data_0_3_7 <= line_write_buffer_data_0[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_312) begin // @[Sbuffer.scala 149:27]
      data_0_3_8 <= line_write_buffer_data_0_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_56) begin // @[Sbuffer.scala 149:27]
      data_0_3_8 <= line_write_buffer_data_0[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_313) begin // @[Sbuffer.scala 149:27]
      data_0_3_9 <= line_write_buffer_data_0_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_57) begin // @[Sbuffer.scala 149:27]
      data_0_3_9 <= line_write_buffer_data_0[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_314) begin // @[Sbuffer.scala 149:27]
      data_0_3_10 <= line_write_buffer_data_0_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_58) begin // @[Sbuffer.scala 149:27]
      data_0_3_10 <= line_write_buffer_data_0[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_315) begin // @[Sbuffer.scala 149:27]
      data_0_3_11 <= line_write_buffer_data_0_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_59) begin // @[Sbuffer.scala 149:27]
      data_0_3_11 <= line_write_buffer_data_0[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_316) begin // @[Sbuffer.scala 149:27]
      data_0_3_12 <= line_write_buffer_data_0_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_60) begin // @[Sbuffer.scala 149:27]
      data_0_3_12 <= line_write_buffer_data_0[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_317) begin // @[Sbuffer.scala 149:27]
      data_0_3_13 <= line_write_buffer_data_0_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_61) begin // @[Sbuffer.scala 149:27]
      data_0_3_13 <= line_write_buffer_data_0[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_318) begin // @[Sbuffer.scala 149:27]
      data_0_3_14 <= line_write_buffer_data_0_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_62) begin // @[Sbuffer.scala 149:27]
      data_0_3_14 <= line_write_buffer_data_0[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_319) begin // @[Sbuffer.scala 149:27]
      data_0_3_15 <= line_write_buffer_data_0_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_63) begin // @[Sbuffer.scala 149:27]
      data_0_3_15 <= line_write_buffer_data_0[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_320) begin // @[Sbuffer.scala 149:27]
      data_1_0_0 <= line_write_buffer_data_1_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_64) begin // @[Sbuffer.scala 149:27]
      data_1_0_0 <= line_write_buffer_data_1[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_321) begin // @[Sbuffer.scala 149:27]
      data_1_0_1 <= line_write_buffer_data_1_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_65) begin // @[Sbuffer.scala 149:27]
      data_1_0_1 <= line_write_buffer_data_1[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_322) begin // @[Sbuffer.scala 149:27]
      data_1_0_2 <= line_write_buffer_data_1_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_66) begin // @[Sbuffer.scala 149:27]
      data_1_0_2 <= line_write_buffer_data_1[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_323) begin // @[Sbuffer.scala 149:27]
      data_1_0_3 <= line_write_buffer_data_1_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_67) begin // @[Sbuffer.scala 149:27]
      data_1_0_3 <= line_write_buffer_data_1[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_324) begin // @[Sbuffer.scala 149:27]
      data_1_0_4 <= line_write_buffer_data_1_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_68) begin // @[Sbuffer.scala 149:27]
      data_1_0_4 <= line_write_buffer_data_1[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_325) begin // @[Sbuffer.scala 149:27]
      data_1_0_5 <= line_write_buffer_data_1_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_69) begin // @[Sbuffer.scala 149:27]
      data_1_0_5 <= line_write_buffer_data_1[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_326) begin // @[Sbuffer.scala 149:27]
      data_1_0_6 <= line_write_buffer_data_1_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_70) begin // @[Sbuffer.scala 149:27]
      data_1_0_6 <= line_write_buffer_data_1[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_327) begin // @[Sbuffer.scala 149:27]
      data_1_0_7 <= line_write_buffer_data_1_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_71) begin // @[Sbuffer.scala 149:27]
      data_1_0_7 <= line_write_buffer_data_1[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_328) begin // @[Sbuffer.scala 149:27]
      data_1_0_8 <= line_write_buffer_data_1_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_72) begin // @[Sbuffer.scala 149:27]
      data_1_0_8 <= line_write_buffer_data_1[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_329) begin // @[Sbuffer.scala 149:27]
      data_1_0_9 <= line_write_buffer_data_1_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_73) begin // @[Sbuffer.scala 149:27]
      data_1_0_9 <= line_write_buffer_data_1[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_330) begin // @[Sbuffer.scala 149:27]
      data_1_0_10 <= line_write_buffer_data_1_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_74) begin // @[Sbuffer.scala 149:27]
      data_1_0_10 <= line_write_buffer_data_1[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_331) begin // @[Sbuffer.scala 149:27]
      data_1_0_11 <= line_write_buffer_data_1_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_75) begin // @[Sbuffer.scala 149:27]
      data_1_0_11 <= line_write_buffer_data_1[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_332) begin // @[Sbuffer.scala 149:27]
      data_1_0_12 <= line_write_buffer_data_1_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_76) begin // @[Sbuffer.scala 149:27]
      data_1_0_12 <= line_write_buffer_data_1[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_333) begin // @[Sbuffer.scala 149:27]
      data_1_0_13 <= line_write_buffer_data_1_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_77) begin // @[Sbuffer.scala 149:27]
      data_1_0_13 <= line_write_buffer_data_1[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_334) begin // @[Sbuffer.scala 149:27]
      data_1_0_14 <= line_write_buffer_data_1_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_78) begin // @[Sbuffer.scala 149:27]
      data_1_0_14 <= line_write_buffer_data_1[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_335) begin // @[Sbuffer.scala 149:27]
      data_1_0_15 <= line_write_buffer_data_1_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_79) begin // @[Sbuffer.scala 149:27]
      data_1_0_15 <= line_write_buffer_data_1[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_336) begin // @[Sbuffer.scala 149:27]
      data_1_1_0 <= line_write_buffer_data_1_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_80) begin // @[Sbuffer.scala 149:27]
      data_1_1_0 <= line_write_buffer_data_1[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_337) begin // @[Sbuffer.scala 149:27]
      data_1_1_1 <= line_write_buffer_data_1_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_81) begin // @[Sbuffer.scala 149:27]
      data_1_1_1 <= line_write_buffer_data_1[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_338) begin // @[Sbuffer.scala 149:27]
      data_1_1_2 <= line_write_buffer_data_1_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_82) begin // @[Sbuffer.scala 149:27]
      data_1_1_2 <= line_write_buffer_data_1[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_339) begin // @[Sbuffer.scala 149:27]
      data_1_1_3 <= line_write_buffer_data_1_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_83) begin // @[Sbuffer.scala 149:27]
      data_1_1_3 <= line_write_buffer_data_1[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_340) begin // @[Sbuffer.scala 149:27]
      data_1_1_4 <= line_write_buffer_data_1_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_84) begin // @[Sbuffer.scala 149:27]
      data_1_1_4 <= line_write_buffer_data_1[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_341) begin // @[Sbuffer.scala 149:27]
      data_1_1_5 <= line_write_buffer_data_1_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_85) begin // @[Sbuffer.scala 149:27]
      data_1_1_5 <= line_write_buffer_data_1[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_342) begin // @[Sbuffer.scala 149:27]
      data_1_1_6 <= line_write_buffer_data_1_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_86) begin // @[Sbuffer.scala 149:27]
      data_1_1_6 <= line_write_buffer_data_1[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_343) begin // @[Sbuffer.scala 149:27]
      data_1_1_7 <= line_write_buffer_data_1_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_87) begin // @[Sbuffer.scala 149:27]
      data_1_1_7 <= line_write_buffer_data_1[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_344) begin // @[Sbuffer.scala 149:27]
      data_1_1_8 <= line_write_buffer_data_1_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_88) begin // @[Sbuffer.scala 149:27]
      data_1_1_8 <= line_write_buffer_data_1[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_345) begin // @[Sbuffer.scala 149:27]
      data_1_1_9 <= line_write_buffer_data_1_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_89) begin // @[Sbuffer.scala 149:27]
      data_1_1_9 <= line_write_buffer_data_1[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_346) begin // @[Sbuffer.scala 149:27]
      data_1_1_10 <= line_write_buffer_data_1_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_90) begin // @[Sbuffer.scala 149:27]
      data_1_1_10 <= line_write_buffer_data_1[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_347) begin // @[Sbuffer.scala 149:27]
      data_1_1_11 <= line_write_buffer_data_1_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_91) begin // @[Sbuffer.scala 149:27]
      data_1_1_11 <= line_write_buffer_data_1[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_348) begin // @[Sbuffer.scala 149:27]
      data_1_1_12 <= line_write_buffer_data_1_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_92) begin // @[Sbuffer.scala 149:27]
      data_1_1_12 <= line_write_buffer_data_1[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_349) begin // @[Sbuffer.scala 149:27]
      data_1_1_13 <= line_write_buffer_data_1_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_93) begin // @[Sbuffer.scala 149:27]
      data_1_1_13 <= line_write_buffer_data_1[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_350) begin // @[Sbuffer.scala 149:27]
      data_1_1_14 <= line_write_buffer_data_1_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_94) begin // @[Sbuffer.scala 149:27]
      data_1_1_14 <= line_write_buffer_data_1[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_351) begin // @[Sbuffer.scala 149:27]
      data_1_1_15 <= line_write_buffer_data_1_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_95) begin // @[Sbuffer.scala 149:27]
      data_1_1_15 <= line_write_buffer_data_1[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_352) begin // @[Sbuffer.scala 149:27]
      data_1_2_0 <= line_write_buffer_data_1_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_96) begin // @[Sbuffer.scala 149:27]
      data_1_2_0 <= line_write_buffer_data_1[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_353) begin // @[Sbuffer.scala 149:27]
      data_1_2_1 <= line_write_buffer_data_1_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_97) begin // @[Sbuffer.scala 149:27]
      data_1_2_1 <= line_write_buffer_data_1[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_354) begin // @[Sbuffer.scala 149:27]
      data_1_2_2 <= line_write_buffer_data_1_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_98) begin // @[Sbuffer.scala 149:27]
      data_1_2_2 <= line_write_buffer_data_1[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_355) begin // @[Sbuffer.scala 149:27]
      data_1_2_3 <= line_write_buffer_data_1_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_99) begin // @[Sbuffer.scala 149:27]
      data_1_2_3 <= line_write_buffer_data_1[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_356) begin // @[Sbuffer.scala 149:27]
      data_1_2_4 <= line_write_buffer_data_1_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_100) begin // @[Sbuffer.scala 149:27]
      data_1_2_4 <= line_write_buffer_data_1[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_357) begin // @[Sbuffer.scala 149:27]
      data_1_2_5 <= line_write_buffer_data_1_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_101) begin // @[Sbuffer.scala 149:27]
      data_1_2_5 <= line_write_buffer_data_1[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_358) begin // @[Sbuffer.scala 149:27]
      data_1_2_6 <= line_write_buffer_data_1_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_102) begin // @[Sbuffer.scala 149:27]
      data_1_2_6 <= line_write_buffer_data_1[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_359) begin // @[Sbuffer.scala 149:27]
      data_1_2_7 <= line_write_buffer_data_1_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_103) begin // @[Sbuffer.scala 149:27]
      data_1_2_7 <= line_write_buffer_data_1[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_360) begin // @[Sbuffer.scala 149:27]
      data_1_2_8 <= line_write_buffer_data_1_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_104) begin // @[Sbuffer.scala 149:27]
      data_1_2_8 <= line_write_buffer_data_1[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_361) begin // @[Sbuffer.scala 149:27]
      data_1_2_9 <= line_write_buffer_data_1_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_105) begin // @[Sbuffer.scala 149:27]
      data_1_2_9 <= line_write_buffer_data_1[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_362) begin // @[Sbuffer.scala 149:27]
      data_1_2_10 <= line_write_buffer_data_1_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_106) begin // @[Sbuffer.scala 149:27]
      data_1_2_10 <= line_write_buffer_data_1[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_363) begin // @[Sbuffer.scala 149:27]
      data_1_2_11 <= line_write_buffer_data_1_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_107) begin // @[Sbuffer.scala 149:27]
      data_1_2_11 <= line_write_buffer_data_1[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_364) begin // @[Sbuffer.scala 149:27]
      data_1_2_12 <= line_write_buffer_data_1_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_108) begin // @[Sbuffer.scala 149:27]
      data_1_2_12 <= line_write_buffer_data_1[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_365) begin // @[Sbuffer.scala 149:27]
      data_1_2_13 <= line_write_buffer_data_1_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_109) begin // @[Sbuffer.scala 149:27]
      data_1_2_13 <= line_write_buffer_data_1[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_366) begin // @[Sbuffer.scala 149:27]
      data_1_2_14 <= line_write_buffer_data_1_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_110) begin // @[Sbuffer.scala 149:27]
      data_1_2_14 <= line_write_buffer_data_1[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_367) begin // @[Sbuffer.scala 149:27]
      data_1_2_15 <= line_write_buffer_data_1_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_111) begin // @[Sbuffer.scala 149:27]
      data_1_2_15 <= line_write_buffer_data_1[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_368) begin // @[Sbuffer.scala 149:27]
      data_1_3_0 <= line_write_buffer_data_1_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_112) begin // @[Sbuffer.scala 149:27]
      data_1_3_0 <= line_write_buffer_data_1[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_369) begin // @[Sbuffer.scala 149:27]
      data_1_3_1 <= line_write_buffer_data_1_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_113) begin // @[Sbuffer.scala 149:27]
      data_1_3_1 <= line_write_buffer_data_1[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_370) begin // @[Sbuffer.scala 149:27]
      data_1_3_2 <= line_write_buffer_data_1_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_114) begin // @[Sbuffer.scala 149:27]
      data_1_3_2 <= line_write_buffer_data_1[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_371) begin // @[Sbuffer.scala 149:27]
      data_1_3_3 <= line_write_buffer_data_1_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_115) begin // @[Sbuffer.scala 149:27]
      data_1_3_3 <= line_write_buffer_data_1[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_372) begin // @[Sbuffer.scala 149:27]
      data_1_3_4 <= line_write_buffer_data_1_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_116) begin // @[Sbuffer.scala 149:27]
      data_1_3_4 <= line_write_buffer_data_1[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_373) begin // @[Sbuffer.scala 149:27]
      data_1_3_5 <= line_write_buffer_data_1_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_117) begin // @[Sbuffer.scala 149:27]
      data_1_3_5 <= line_write_buffer_data_1[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_374) begin // @[Sbuffer.scala 149:27]
      data_1_3_6 <= line_write_buffer_data_1_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_118) begin // @[Sbuffer.scala 149:27]
      data_1_3_6 <= line_write_buffer_data_1[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_375) begin // @[Sbuffer.scala 149:27]
      data_1_3_7 <= line_write_buffer_data_1_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_119) begin // @[Sbuffer.scala 149:27]
      data_1_3_7 <= line_write_buffer_data_1[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_376) begin // @[Sbuffer.scala 149:27]
      data_1_3_8 <= line_write_buffer_data_1_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_120) begin // @[Sbuffer.scala 149:27]
      data_1_3_8 <= line_write_buffer_data_1[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_377) begin // @[Sbuffer.scala 149:27]
      data_1_3_9 <= line_write_buffer_data_1_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_121) begin // @[Sbuffer.scala 149:27]
      data_1_3_9 <= line_write_buffer_data_1[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_378) begin // @[Sbuffer.scala 149:27]
      data_1_3_10 <= line_write_buffer_data_1_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_122) begin // @[Sbuffer.scala 149:27]
      data_1_3_10 <= line_write_buffer_data_1[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_379) begin // @[Sbuffer.scala 149:27]
      data_1_3_11 <= line_write_buffer_data_1_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_123) begin // @[Sbuffer.scala 149:27]
      data_1_3_11 <= line_write_buffer_data_1[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_380) begin // @[Sbuffer.scala 149:27]
      data_1_3_12 <= line_write_buffer_data_1_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_124) begin // @[Sbuffer.scala 149:27]
      data_1_3_12 <= line_write_buffer_data_1[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_381) begin // @[Sbuffer.scala 149:27]
      data_1_3_13 <= line_write_buffer_data_1_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_125) begin // @[Sbuffer.scala 149:27]
      data_1_3_13 <= line_write_buffer_data_1[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_382) begin // @[Sbuffer.scala 149:27]
      data_1_3_14 <= line_write_buffer_data_1_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_126) begin // @[Sbuffer.scala 149:27]
      data_1_3_14 <= line_write_buffer_data_1[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_383) begin // @[Sbuffer.scala 149:27]
      data_1_3_15 <= line_write_buffer_data_1_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_127) begin // @[Sbuffer.scala 149:27]
      data_1_3_15 <= line_write_buffer_data_1[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_384) begin // @[Sbuffer.scala 149:27]
      data_2_0_0 <= line_write_buffer_data_2_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_128) begin // @[Sbuffer.scala 149:27]
      data_2_0_0 <= line_write_buffer_data_2[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_385) begin // @[Sbuffer.scala 149:27]
      data_2_0_1 <= line_write_buffer_data_2_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_129) begin // @[Sbuffer.scala 149:27]
      data_2_0_1 <= line_write_buffer_data_2[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_386) begin // @[Sbuffer.scala 149:27]
      data_2_0_2 <= line_write_buffer_data_2_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_130) begin // @[Sbuffer.scala 149:27]
      data_2_0_2 <= line_write_buffer_data_2[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_387) begin // @[Sbuffer.scala 149:27]
      data_2_0_3 <= line_write_buffer_data_2_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_131) begin // @[Sbuffer.scala 149:27]
      data_2_0_3 <= line_write_buffer_data_2[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_388) begin // @[Sbuffer.scala 149:27]
      data_2_0_4 <= line_write_buffer_data_2_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_132) begin // @[Sbuffer.scala 149:27]
      data_2_0_4 <= line_write_buffer_data_2[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_389) begin // @[Sbuffer.scala 149:27]
      data_2_0_5 <= line_write_buffer_data_2_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_133) begin // @[Sbuffer.scala 149:27]
      data_2_0_5 <= line_write_buffer_data_2[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_390) begin // @[Sbuffer.scala 149:27]
      data_2_0_6 <= line_write_buffer_data_2_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_134) begin // @[Sbuffer.scala 149:27]
      data_2_0_6 <= line_write_buffer_data_2[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_391) begin // @[Sbuffer.scala 149:27]
      data_2_0_7 <= line_write_buffer_data_2_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_135) begin // @[Sbuffer.scala 149:27]
      data_2_0_7 <= line_write_buffer_data_2[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_392) begin // @[Sbuffer.scala 149:27]
      data_2_0_8 <= line_write_buffer_data_2_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_136) begin // @[Sbuffer.scala 149:27]
      data_2_0_8 <= line_write_buffer_data_2[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_393) begin // @[Sbuffer.scala 149:27]
      data_2_0_9 <= line_write_buffer_data_2_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_137) begin // @[Sbuffer.scala 149:27]
      data_2_0_9 <= line_write_buffer_data_2[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_394) begin // @[Sbuffer.scala 149:27]
      data_2_0_10 <= line_write_buffer_data_2_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_138) begin // @[Sbuffer.scala 149:27]
      data_2_0_10 <= line_write_buffer_data_2[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_395) begin // @[Sbuffer.scala 149:27]
      data_2_0_11 <= line_write_buffer_data_2_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_139) begin // @[Sbuffer.scala 149:27]
      data_2_0_11 <= line_write_buffer_data_2[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_396) begin // @[Sbuffer.scala 149:27]
      data_2_0_12 <= line_write_buffer_data_2_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_140) begin // @[Sbuffer.scala 149:27]
      data_2_0_12 <= line_write_buffer_data_2[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_397) begin // @[Sbuffer.scala 149:27]
      data_2_0_13 <= line_write_buffer_data_2_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_141) begin // @[Sbuffer.scala 149:27]
      data_2_0_13 <= line_write_buffer_data_2[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_398) begin // @[Sbuffer.scala 149:27]
      data_2_0_14 <= line_write_buffer_data_2_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_142) begin // @[Sbuffer.scala 149:27]
      data_2_0_14 <= line_write_buffer_data_2[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_399) begin // @[Sbuffer.scala 149:27]
      data_2_0_15 <= line_write_buffer_data_2_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_143) begin // @[Sbuffer.scala 149:27]
      data_2_0_15 <= line_write_buffer_data_2[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_400) begin // @[Sbuffer.scala 149:27]
      data_2_1_0 <= line_write_buffer_data_2_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_144) begin // @[Sbuffer.scala 149:27]
      data_2_1_0 <= line_write_buffer_data_2[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_401) begin // @[Sbuffer.scala 149:27]
      data_2_1_1 <= line_write_buffer_data_2_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_145) begin // @[Sbuffer.scala 149:27]
      data_2_1_1 <= line_write_buffer_data_2[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_402) begin // @[Sbuffer.scala 149:27]
      data_2_1_2 <= line_write_buffer_data_2_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_146) begin // @[Sbuffer.scala 149:27]
      data_2_1_2 <= line_write_buffer_data_2[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_403) begin // @[Sbuffer.scala 149:27]
      data_2_1_3 <= line_write_buffer_data_2_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_147) begin // @[Sbuffer.scala 149:27]
      data_2_1_3 <= line_write_buffer_data_2[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_404) begin // @[Sbuffer.scala 149:27]
      data_2_1_4 <= line_write_buffer_data_2_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_148) begin // @[Sbuffer.scala 149:27]
      data_2_1_4 <= line_write_buffer_data_2[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_405) begin // @[Sbuffer.scala 149:27]
      data_2_1_5 <= line_write_buffer_data_2_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_149) begin // @[Sbuffer.scala 149:27]
      data_2_1_5 <= line_write_buffer_data_2[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_406) begin // @[Sbuffer.scala 149:27]
      data_2_1_6 <= line_write_buffer_data_2_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_150) begin // @[Sbuffer.scala 149:27]
      data_2_1_6 <= line_write_buffer_data_2[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_407) begin // @[Sbuffer.scala 149:27]
      data_2_1_7 <= line_write_buffer_data_2_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_151) begin // @[Sbuffer.scala 149:27]
      data_2_1_7 <= line_write_buffer_data_2[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_408) begin // @[Sbuffer.scala 149:27]
      data_2_1_8 <= line_write_buffer_data_2_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_152) begin // @[Sbuffer.scala 149:27]
      data_2_1_8 <= line_write_buffer_data_2[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_409) begin // @[Sbuffer.scala 149:27]
      data_2_1_9 <= line_write_buffer_data_2_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_153) begin // @[Sbuffer.scala 149:27]
      data_2_1_9 <= line_write_buffer_data_2[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_410) begin // @[Sbuffer.scala 149:27]
      data_2_1_10 <= line_write_buffer_data_2_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_154) begin // @[Sbuffer.scala 149:27]
      data_2_1_10 <= line_write_buffer_data_2[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_411) begin // @[Sbuffer.scala 149:27]
      data_2_1_11 <= line_write_buffer_data_2_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_155) begin // @[Sbuffer.scala 149:27]
      data_2_1_11 <= line_write_buffer_data_2[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_412) begin // @[Sbuffer.scala 149:27]
      data_2_1_12 <= line_write_buffer_data_2_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_156) begin // @[Sbuffer.scala 149:27]
      data_2_1_12 <= line_write_buffer_data_2[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_413) begin // @[Sbuffer.scala 149:27]
      data_2_1_13 <= line_write_buffer_data_2_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_157) begin // @[Sbuffer.scala 149:27]
      data_2_1_13 <= line_write_buffer_data_2[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_414) begin // @[Sbuffer.scala 149:27]
      data_2_1_14 <= line_write_buffer_data_2_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_158) begin // @[Sbuffer.scala 149:27]
      data_2_1_14 <= line_write_buffer_data_2[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_415) begin // @[Sbuffer.scala 149:27]
      data_2_1_15 <= line_write_buffer_data_2_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_159) begin // @[Sbuffer.scala 149:27]
      data_2_1_15 <= line_write_buffer_data_2[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_416) begin // @[Sbuffer.scala 149:27]
      data_2_2_0 <= line_write_buffer_data_2_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_160) begin // @[Sbuffer.scala 149:27]
      data_2_2_0 <= line_write_buffer_data_2[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_417) begin // @[Sbuffer.scala 149:27]
      data_2_2_1 <= line_write_buffer_data_2_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_161) begin // @[Sbuffer.scala 149:27]
      data_2_2_1 <= line_write_buffer_data_2[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_418) begin // @[Sbuffer.scala 149:27]
      data_2_2_2 <= line_write_buffer_data_2_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_162) begin // @[Sbuffer.scala 149:27]
      data_2_2_2 <= line_write_buffer_data_2[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_419) begin // @[Sbuffer.scala 149:27]
      data_2_2_3 <= line_write_buffer_data_2_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_163) begin // @[Sbuffer.scala 149:27]
      data_2_2_3 <= line_write_buffer_data_2[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_420) begin // @[Sbuffer.scala 149:27]
      data_2_2_4 <= line_write_buffer_data_2_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_164) begin // @[Sbuffer.scala 149:27]
      data_2_2_4 <= line_write_buffer_data_2[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_421) begin // @[Sbuffer.scala 149:27]
      data_2_2_5 <= line_write_buffer_data_2_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_165) begin // @[Sbuffer.scala 149:27]
      data_2_2_5 <= line_write_buffer_data_2[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_422) begin // @[Sbuffer.scala 149:27]
      data_2_2_6 <= line_write_buffer_data_2_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_166) begin // @[Sbuffer.scala 149:27]
      data_2_2_6 <= line_write_buffer_data_2[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_423) begin // @[Sbuffer.scala 149:27]
      data_2_2_7 <= line_write_buffer_data_2_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_167) begin // @[Sbuffer.scala 149:27]
      data_2_2_7 <= line_write_buffer_data_2[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_424) begin // @[Sbuffer.scala 149:27]
      data_2_2_8 <= line_write_buffer_data_2_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_168) begin // @[Sbuffer.scala 149:27]
      data_2_2_8 <= line_write_buffer_data_2[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_425) begin // @[Sbuffer.scala 149:27]
      data_2_2_9 <= line_write_buffer_data_2_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_169) begin // @[Sbuffer.scala 149:27]
      data_2_2_9 <= line_write_buffer_data_2[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_426) begin // @[Sbuffer.scala 149:27]
      data_2_2_10 <= line_write_buffer_data_2_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_170) begin // @[Sbuffer.scala 149:27]
      data_2_2_10 <= line_write_buffer_data_2[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_427) begin // @[Sbuffer.scala 149:27]
      data_2_2_11 <= line_write_buffer_data_2_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_171) begin // @[Sbuffer.scala 149:27]
      data_2_2_11 <= line_write_buffer_data_2[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_428) begin // @[Sbuffer.scala 149:27]
      data_2_2_12 <= line_write_buffer_data_2_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_172) begin // @[Sbuffer.scala 149:27]
      data_2_2_12 <= line_write_buffer_data_2[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_429) begin // @[Sbuffer.scala 149:27]
      data_2_2_13 <= line_write_buffer_data_2_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_173) begin // @[Sbuffer.scala 149:27]
      data_2_2_13 <= line_write_buffer_data_2[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_430) begin // @[Sbuffer.scala 149:27]
      data_2_2_14 <= line_write_buffer_data_2_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_174) begin // @[Sbuffer.scala 149:27]
      data_2_2_14 <= line_write_buffer_data_2[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_431) begin // @[Sbuffer.scala 149:27]
      data_2_2_15 <= line_write_buffer_data_2_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_175) begin // @[Sbuffer.scala 149:27]
      data_2_2_15 <= line_write_buffer_data_2[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_432) begin // @[Sbuffer.scala 149:27]
      data_2_3_0 <= line_write_buffer_data_2_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_176) begin // @[Sbuffer.scala 149:27]
      data_2_3_0 <= line_write_buffer_data_2[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_433) begin // @[Sbuffer.scala 149:27]
      data_2_3_1 <= line_write_buffer_data_2_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_177) begin // @[Sbuffer.scala 149:27]
      data_2_3_1 <= line_write_buffer_data_2[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_434) begin // @[Sbuffer.scala 149:27]
      data_2_3_2 <= line_write_buffer_data_2_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_178) begin // @[Sbuffer.scala 149:27]
      data_2_3_2 <= line_write_buffer_data_2[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_435) begin // @[Sbuffer.scala 149:27]
      data_2_3_3 <= line_write_buffer_data_2_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_179) begin // @[Sbuffer.scala 149:27]
      data_2_3_3 <= line_write_buffer_data_2[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_436) begin // @[Sbuffer.scala 149:27]
      data_2_3_4 <= line_write_buffer_data_2_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_180) begin // @[Sbuffer.scala 149:27]
      data_2_3_4 <= line_write_buffer_data_2[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_437) begin // @[Sbuffer.scala 149:27]
      data_2_3_5 <= line_write_buffer_data_2_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_181) begin // @[Sbuffer.scala 149:27]
      data_2_3_5 <= line_write_buffer_data_2[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_438) begin // @[Sbuffer.scala 149:27]
      data_2_3_6 <= line_write_buffer_data_2_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_182) begin // @[Sbuffer.scala 149:27]
      data_2_3_6 <= line_write_buffer_data_2[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_439) begin // @[Sbuffer.scala 149:27]
      data_2_3_7 <= line_write_buffer_data_2_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_183) begin // @[Sbuffer.scala 149:27]
      data_2_3_7 <= line_write_buffer_data_2[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_440) begin // @[Sbuffer.scala 149:27]
      data_2_3_8 <= line_write_buffer_data_2_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_184) begin // @[Sbuffer.scala 149:27]
      data_2_3_8 <= line_write_buffer_data_2[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_441) begin // @[Sbuffer.scala 149:27]
      data_2_3_9 <= line_write_buffer_data_2_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_185) begin // @[Sbuffer.scala 149:27]
      data_2_3_9 <= line_write_buffer_data_2[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_442) begin // @[Sbuffer.scala 149:27]
      data_2_3_10 <= line_write_buffer_data_2_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_186) begin // @[Sbuffer.scala 149:27]
      data_2_3_10 <= line_write_buffer_data_2[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_443) begin // @[Sbuffer.scala 149:27]
      data_2_3_11 <= line_write_buffer_data_2_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_187) begin // @[Sbuffer.scala 149:27]
      data_2_3_11 <= line_write_buffer_data_2[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_444) begin // @[Sbuffer.scala 149:27]
      data_2_3_12 <= line_write_buffer_data_2_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_188) begin // @[Sbuffer.scala 149:27]
      data_2_3_12 <= line_write_buffer_data_2[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_445) begin // @[Sbuffer.scala 149:27]
      data_2_3_13 <= line_write_buffer_data_2_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_189) begin // @[Sbuffer.scala 149:27]
      data_2_3_13 <= line_write_buffer_data_2[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_446) begin // @[Sbuffer.scala 149:27]
      data_2_3_14 <= line_write_buffer_data_2_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_190) begin // @[Sbuffer.scala 149:27]
      data_2_3_14 <= line_write_buffer_data_2[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_447) begin // @[Sbuffer.scala 149:27]
      data_2_3_15 <= line_write_buffer_data_2_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_191) begin // @[Sbuffer.scala 149:27]
      data_2_3_15 <= line_write_buffer_data_2[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_448) begin // @[Sbuffer.scala 149:27]
      data_3_0_0 <= line_write_buffer_data_3_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_192) begin // @[Sbuffer.scala 149:27]
      data_3_0_0 <= line_write_buffer_data_3[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_449) begin // @[Sbuffer.scala 149:27]
      data_3_0_1 <= line_write_buffer_data_3_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_193) begin // @[Sbuffer.scala 149:27]
      data_3_0_1 <= line_write_buffer_data_3[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_450) begin // @[Sbuffer.scala 149:27]
      data_3_0_2 <= line_write_buffer_data_3_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_194) begin // @[Sbuffer.scala 149:27]
      data_3_0_2 <= line_write_buffer_data_3[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_451) begin // @[Sbuffer.scala 149:27]
      data_3_0_3 <= line_write_buffer_data_3_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_195) begin // @[Sbuffer.scala 149:27]
      data_3_0_3 <= line_write_buffer_data_3[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_452) begin // @[Sbuffer.scala 149:27]
      data_3_0_4 <= line_write_buffer_data_3_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_196) begin // @[Sbuffer.scala 149:27]
      data_3_0_4 <= line_write_buffer_data_3[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_453) begin // @[Sbuffer.scala 149:27]
      data_3_0_5 <= line_write_buffer_data_3_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_197) begin // @[Sbuffer.scala 149:27]
      data_3_0_5 <= line_write_buffer_data_3[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_454) begin // @[Sbuffer.scala 149:27]
      data_3_0_6 <= line_write_buffer_data_3_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_198) begin // @[Sbuffer.scala 149:27]
      data_3_0_6 <= line_write_buffer_data_3[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_455) begin // @[Sbuffer.scala 149:27]
      data_3_0_7 <= line_write_buffer_data_3_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_199) begin // @[Sbuffer.scala 149:27]
      data_3_0_7 <= line_write_buffer_data_3[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_456) begin // @[Sbuffer.scala 149:27]
      data_3_0_8 <= line_write_buffer_data_3_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_200) begin // @[Sbuffer.scala 149:27]
      data_3_0_8 <= line_write_buffer_data_3[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_457) begin // @[Sbuffer.scala 149:27]
      data_3_0_9 <= line_write_buffer_data_3_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_201) begin // @[Sbuffer.scala 149:27]
      data_3_0_9 <= line_write_buffer_data_3[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_458) begin // @[Sbuffer.scala 149:27]
      data_3_0_10 <= line_write_buffer_data_3_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_202) begin // @[Sbuffer.scala 149:27]
      data_3_0_10 <= line_write_buffer_data_3[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_459) begin // @[Sbuffer.scala 149:27]
      data_3_0_11 <= line_write_buffer_data_3_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_203) begin // @[Sbuffer.scala 149:27]
      data_3_0_11 <= line_write_buffer_data_3[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_460) begin // @[Sbuffer.scala 149:27]
      data_3_0_12 <= line_write_buffer_data_3_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_204) begin // @[Sbuffer.scala 149:27]
      data_3_0_12 <= line_write_buffer_data_3[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_461) begin // @[Sbuffer.scala 149:27]
      data_3_0_13 <= line_write_buffer_data_3_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_205) begin // @[Sbuffer.scala 149:27]
      data_3_0_13 <= line_write_buffer_data_3[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_462) begin // @[Sbuffer.scala 149:27]
      data_3_0_14 <= line_write_buffer_data_3_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_206) begin // @[Sbuffer.scala 149:27]
      data_3_0_14 <= line_write_buffer_data_3[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_463) begin // @[Sbuffer.scala 149:27]
      data_3_0_15 <= line_write_buffer_data_3_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_207) begin // @[Sbuffer.scala 149:27]
      data_3_0_15 <= line_write_buffer_data_3[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_464) begin // @[Sbuffer.scala 149:27]
      data_3_1_0 <= line_write_buffer_data_3_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_208) begin // @[Sbuffer.scala 149:27]
      data_3_1_0 <= line_write_buffer_data_3[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_465) begin // @[Sbuffer.scala 149:27]
      data_3_1_1 <= line_write_buffer_data_3_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_209) begin // @[Sbuffer.scala 149:27]
      data_3_1_1 <= line_write_buffer_data_3[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_466) begin // @[Sbuffer.scala 149:27]
      data_3_1_2 <= line_write_buffer_data_3_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_210) begin // @[Sbuffer.scala 149:27]
      data_3_1_2 <= line_write_buffer_data_3[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_467) begin // @[Sbuffer.scala 149:27]
      data_3_1_3 <= line_write_buffer_data_3_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_211) begin // @[Sbuffer.scala 149:27]
      data_3_1_3 <= line_write_buffer_data_3[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_468) begin // @[Sbuffer.scala 149:27]
      data_3_1_4 <= line_write_buffer_data_3_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_212) begin // @[Sbuffer.scala 149:27]
      data_3_1_4 <= line_write_buffer_data_3[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_469) begin // @[Sbuffer.scala 149:27]
      data_3_1_5 <= line_write_buffer_data_3_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_213) begin // @[Sbuffer.scala 149:27]
      data_3_1_5 <= line_write_buffer_data_3[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_470) begin // @[Sbuffer.scala 149:27]
      data_3_1_6 <= line_write_buffer_data_3_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_214) begin // @[Sbuffer.scala 149:27]
      data_3_1_6 <= line_write_buffer_data_3[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_471) begin // @[Sbuffer.scala 149:27]
      data_3_1_7 <= line_write_buffer_data_3_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_215) begin // @[Sbuffer.scala 149:27]
      data_3_1_7 <= line_write_buffer_data_3[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_472) begin // @[Sbuffer.scala 149:27]
      data_3_1_8 <= line_write_buffer_data_3_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_216) begin // @[Sbuffer.scala 149:27]
      data_3_1_8 <= line_write_buffer_data_3[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_473) begin // @[Sbuffer.scala 149:27]
      data_3_1_9 <= line_write_buffer_data_3_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_217) begin // @[Sbuffer.scala 149:27]
      data_3_1_9 <= line_write_buffer_data_3[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_474) begin // @[Sbuffer.scala 149:27]
      data_3_1_10 <= line_write_buffer_data_3_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_218) begin // @[Sbuffer.scala 149:27]
      data_3_1_10 <= line_write_buffer_data_3[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_475) begin // @[Sbuffer.scala 149:27]
      data_3_1_11 <= line_write_buffer_data_3_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_219) begin // @[Sbuffer.scala 149:27]
      data_3_1_11 <= line_write_buffer_data_3[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_476) begin // @[Sbuffer.scala 149:27]
      data_3_1_12 <= line_write_buffer_data_3_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_220) begin // @[Sbuffer.scala 149:27]
      data_3_1_12 <= line_write_buffer_data_3[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_477) begin // @[Sbuffer.scala 149:27]
      data_3_1_13 <= line_write_buffer_data_3_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_221) begin // @[Sbuffer.scala 149:27]
      data_3_1_13 <= line_write_buffer_data_3[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_478) begin // @[Sbuffer.scala 149:27]
      data_3_1_14 <= line_write_buffer_data_3_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_222) begin // @[Sbuffer.scala 149:27]
      data_3_1_14 <= line_write_buffer_data_3[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_479) begin // @[Sbuffer.scala 149:27]
      data_3_1_15 <= line_write_buffer_data_3_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_223) begin // @[Sbuffer.scala 149:27]
      data_3_1_15 <= line_write_buffer_data_3[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_480) begin // @[Sbuffer.scala 149:27]
      data_3_2_0 <= line_write_buffer_data_3_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_224) begin // @[Sbuffer.scala 149:27]
      data_3_2_0 <= line_write_buffer_data_3[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_481) begin // @[Sbuffer.scala 149:27]
      data_3_2_1 <= line_write_buffer_data_3_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_225) begin // @[Sbuffer.scala 149:27]
      data_3_2_1 <= line_write_buffer_data_3[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_482) begin // @[Sbuffer.scala 149:27]
      data_3_2_2 <= line_write_buffer_data_3_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_226) begin // @[Sbuffer.scala 149:27]
      data_3_2_2 <= line_write_buffer_data_3[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_483) begin // @[Sbuffer.scala 149:27]
      data_3_2_3 <= line_write_buffer_data_3_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_227) begin // @[Sbuffer.scala 149:27]
      data_3_2_3 <= line_write_buffer_data_3[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_484) begin // @[Sbuffer.scala 149:27]
      data_3_2_4 <= line_write_buffer_data_3_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_228) begin // @[Sbuffer.scala 149:27]
      data_3_2_4 <= line_write_buffer_data_3[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_485) begin // @[Sbuffer.scala 149:27]
      data_3_2_5 <= line_write_buffer_data_3_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_229) begin // @[Sbuffer.scala 149:27]
      data_3_2_5 <= line_write_buffer_data_3[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_486) begin // @[Sbuffer.scala 149:27]
      data_3_2_6 <= line_write_buffer_data_3_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_230) begin // @[Sbuffer.scala 149:27]
      data_3_2_6 <= line_write_buffer_data_3[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_487) begin // @[Sbuffer.scala 149:27]
      data_3_2_7 <= line_write_buffer_data_3_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_231) begin // @[Sbuffer.scala 149:27]
      data_3_2_7 <= line_write_buffer_data_3[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_488) begin // @[Sbuffer.scala 149:27]
      data_3_2_8 <= line_write_buffer_data_3_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_232) begin // @[Sbuffer.scala 149:27]
      data_3_2_8 <= line_write_buffer_data_3[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_489) begin // @[Sbuffer.scala 149:27]
      data_3_2_9 <= line_write_buffer_data_3_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_233) begin // @[Sbuffer.scala 149:27]
      data_3_2_9 <= line_write_buffer_data_3[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_490) begin // @[Sbuffer.scala 149:27]
      data_3_2_10 <= line_write_buffer_data_3_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_234) begin // @[Sbuffer.scala 149:27]
      data_3_2_10 <= line_write_buffer_data_3[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_491) begin // @[Sbuffer.scala 149:27]
      data_3_2_11 <= line_write_buffer_data_3_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_235) begin // @[Sbuffer.scala 149:27]
      data_3_2_11 <= line_write_buffer_data_3[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_492) begin // @[Sbuffer.scala 149:27]
      data_3_2_12 <= line_write_buffer_data_3_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_236) begin // @[Sbuffer.scala 149:27]
      data_3_2_12 <= line_write_buffer_data_3[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_493) begin // @[Sbuffer.scala 149:27]
      data_3_2_13 <= line_write_buffer_data_3_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_237) begin // @[Sbuffer.scala 149:27]
      data_3_2_13 <= line_write_buffer_data_3[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_494) begin // @[Sbuffer.scala 149:27]
      data_3_2_14 <= line_write_buffer_data_3_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_238) begin // @[Sbuffer.scala 149:27]
      data_3_2_14 <= line_write_buffer_data_3[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_495) begin // @[Sbuffer.scala 149:27]
      data_3_2_15 <= line_write_buffer_data_3_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_239) begin // @[Sbuffer.scala 149:27]
      data_3_2_15 <= line_write_buffer_data_3[127:120]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_496) begin // @[Sbuffer.scala 149:27]
      data_3_3_0 <= line_write_buffer_data_3_1[7:0]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_240) begin // @[Sbuffer.scala 149:27]
      data_3_3_0 <= line_write_buffer_data_3[7:0]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_497) begin // @[Sbuffer.scala 149:27]
      data_3_3_1 <= line_write_buffer_data_3_1[15:8]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_241) begin // @[Sbuffer.scala 149:27]
      data_3_3_1 <= line_write_buffer_data_3[15:8]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_498) begin // @[Sbuffer.scala 149:27]
      data_3_3_2 <= line_write_buffer_data_3_1[23:16]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_242) begin // @[Sbuffer.scala 149:27]
      data_3_3_2 <= line_write_buffer_data_3[23:16]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_499) begin // @[Sbuffer.scala 149:27]
      data_3_3_3 <= line_write_buffer_data_3_1[31:24]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_243) begin // @[Sbuffer.scala 149:27]
      data_3_3_3 <= line_write_buffer_data_3[31:24]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_500) begin // @[Sbuffer.scala 149:27]
      data_3_3_4 <= line_write_buffer_data_3_1[39:32]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_244) begin // @[Sbuffer.scala 149:27]
      data_3_3_4 <= line_write_buffer_data_3[39:32]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_501) begin // @[Sbuffer.scala 149:27]
      data_3_3_5 <= line_write_buffer_data_3_1[47:40]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_245) begin // @[Sbuffer.scala 149:27]
      data_3_3_5 <= line_write_buffer_data_3[47:40]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_502) begin // @[Sbuffer.scala 149:27]
      data_3_3_6 <= line_write_buffer_data_3_1[55:48]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_246) begin // @[Sbuffer.scala 149:27]
      data_3_3_6 <= line_write_buffer_data_3[55:48]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_503) begin // @[Sbuffer.scala 149:27]
      data_3_3_7 <= line_write_buffer_data_3_1[63:56]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_247) begin // @[Sbuffer.scala 149:27]
      data_3_3_7 <= line_write_buffer_data_3[63:56]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_504) begin // @[Sbuffer.scala 149:27]
      data_3_3_8 <= line_write_buffer_data_3_1[71:64]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_248) begin // @[Sbuffer.scala 149:27]
      data_3_3_8 <= line_write_buffer_data_3[71:64]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_505) begin // @[Sbuffer.scala 149:27]
      data_3_3_9 <= line_write_buffer_data_3_1[79:72]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_249) begin // @[Sbuffer.scala 149:27]
      data_3_3_9 <= line_write_buffer_data_3[79:72]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_506) begin // @[Sbuffer.scala 149:27]
      data_3_3_10 <= line_write_buffer_data_3_1[87:80]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_250) begin // @[Sbuffer.scala 149:27]
      data_3_3_10 <= line_write_buffer_data_3[87:80]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_507) begin // @[Sbuffer.scala 149:27]
      data_3_3_11 <= line_write_buffer_data_3_1[95:88]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_251) begin // @[Sbuffer.scala 149:27]
      data_3_3_11 <= line_write_buffer_data_3[95:88]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_508) begin // @[Sbuffer.scala 149:27]
      data_3_3_12 <= line_write_buffer_data_3_1[103:96]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_252) begin // @[Sbuffer.scala 149:27]
      data_3_3_12 <= line_write_buffer_data_3[103:96]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_509) begin // @[Sbuffer.scala 149:27]
      data_3_3_13 <= line_write_buffer_data_3_1[111:104]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_253) begin // @[Sbuffer.scala 149:27]
      data_3_3_13 <= line_write_buffer_data_3[111:104]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_510) begin // @[Sbuffer.scala 149:27]
      data_3_3_14 <= line_write_buffer_data_3_1[119:112]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_254) begin // @[Sbuffer.scala 149:27]
      data_3_3_14 <= line_write_buffer_data_3[119:112]; // @[Sbuffer.scala 150:36]
    end
    if (write_byte_511) begin // @[Sbuffer.scala 149:27]
      data_3_3_15 <= line_write_buffer_data_3_1[127:120]; // @[Sbuffer.scala 150:36]
    end else if (write_byte_255) begin // @[Sbuffer.scala 149:27]
      data_3_3_15 <= line_write_buffer_data_3[127:120]; // @[Sbuffer.scala 150:36]
    end
    line_mask_clean_flag_0 <= io_maskFlushReq_0_valid & io_maskFlushReq_0_bits_wvec[0] | io_maskFlushReq_1_valid &
      io_maskFlushReq_1_bits_wvec[0]; // @[Sbuffer.scala 115:71]
    line_mask_clean_flag_1 <= io_maskFlushReq_0_valid & io_maskFlushReq_0_bits_wvec[1] | io_maskFlushReq_1_valid &
      io_maskFlushReq_1_bits_wvec[1]; // @[Sbuffer.scala 115:71]
    line_mask_clean_flag_2 <= io_maskFlushReq_0_valid & io_maskFlushReq_0_bits_wvec[2] | io_maskFlushReq_1_valid &
      io_maskFlushReq_1_bits_wvec[2]; // @[Sbuffer.scala 115:71]
    line_mask_clean_flag_3 <= io_maskFlushReq_0_valid & io_maskFlushReq_0_bits_wvec[3] | io_maskFlushReq_1_valid &
      io_maskFlushReq_1_bits_wvec[3]; // @[Sbuffer.scala 115:71]
    sbuffer_in_s2_line_wen_0 <= io_writeReq_0_valid & io_writeReq_0_bits_wvec[0]; // @[Sbuffer.scala 131:46]
    if (sbuffer_in_s1_line_wen_0) begin // @[Reg.scala 17:18]
      line_write_buffer_data_0 <= io_writeReq_0_bits_data; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_0) begin // @[Reg.scala 17:18]
      line_write_buffer_wline_0 <= io_writeReq_0_bits_wline; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_0) begin // @[Reg.scala 17:18]
      line_write_buffer_mask_0 <= io_writeReq_0_bits_mask; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_0) begin // @[Reg.scala 17:18]
      line_write_buffer_offset_0 <= io_writeReq_0_bits_vwordOffset[1:0]; // @[Reg.scala 17:22]
    end
    sbuffer_in_s2_line_wen_1 <= io_writeReq_0_valid & io_writeReq_0_bits_wvec[1]; // @[Sbuffer.scala 131:46]
    if (sbuffer_in_s1_line_wen_1) begin // @[Reg.scala 17:18]
      line_write_buffer_data_1 <= io_writeReq_0_bits_data; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_1) begin // @[Reg.scala 17:18]
      line_write_buffer_wline_1 <= io_writeReq_0_bits_wline; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_1) begin // @[Reg.scala 17:18]
      line_write_buffer_mask_1 <= io_writeReq_0_bits_mask; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_1) begin // @[Reg.scala 17:18]
      line_write_buffer_offset_1 <= io_writeReq_0_bits_vwordOffset[1:0]; // @[Reg.scala 17:22]
    end
    sbuffer_in_s2_line_wen_2 <= io_writeReq_0_valid & io_writeReq_0_bits_wvec[2]; // @[Sbuffer.scala 131:46]
    if (sbuffer_in_s1_line_wen_2) begin // @[Reg.scala 17:18]
      line_write_buffer_data_2 <= io_writeReq_0_bits_data; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_2) begin // @[Reg.scala 17:18]
      line_write_buffer_wline_2 <= io_writeReq_0_bits_wline; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_2) begin // @[Reg.scala 17:18]
      line_write_buffer_mask_2 <= io_writeReq_0_bits_mask; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_2) begin // @[Reg.scala 17:18]
      line_write_buffer_offset_2 <= io_writeReq_0_bits_vwordOffset[1:0]; // @[Reg.scala 17:22]
    end
    sbuffer_in_s2_line_wen_3 <= io_writeReq_0_valid & io_writeReq_0_bits_wvec[3]; // @[Sbuffer.scala 131:46]
    if (sbuffer_in_s1_line_wen_3) begin // @[Reg.scala 17:18]
      line_write_buffer_data_3 <= io_writeReq_0_bits_data; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_3) begin // @[Reg.scala 17:18]
      line_write_buffer_wline_3 <= io_writeReq_0_bits_wline; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_3) begin // @[Reg.scala 17:18]
      line_write_buffer_mask_3 <= io_writeReq_0_bits_mask; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_3) begin // @[Reg.scala 17:18]
      line_write_buffer_offset_3 <= io_writeReq_0_bits_vwordOffset[1:0]; // @[Reg.scala 17:22]
    end
    sbuffer_in_s2_line_wen_0_1 <= io_writeReq_1_valid & io_writeReq_1_bits_wvec[0]; // @[Sbuffer.scala 131:46]
    if (sbuffer_in_s1_line_wen_0_1) begin // @[Reg.scala 17:18]
      line_write_buffer_data_0_1 <= io_writeReq_1_bits_data; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_0_1) begin // @[Reg.scala 17:18]
      line_write_buffer_wline_0_1 <= io_writeReq_1_bits_wline; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_0_1) begin // @[Reg.scala 17:18]
      line_write_buffer_mask_0_1 <= io_writeReq_1_bits_mask; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_0_1) begin // @[Reg.scala 17:18]
      line_write_buffer_offset_0_1 <= io_writeReq_1_bits_vwordOffset[1:0]; // @[Reg.scala 17:22]
    end
    sbuffer_in_s2_line_wen_1_1 <= io_writeReq_1_valid & io_writeReq_1_bits_wvec[1]; // @[Sbuffer.scala 131:46]
    if (sbuffer_in_s1_line_wen_1_1) begin // @[Reg.scala 17:18]
      line_write_buffer_data_1_1 <= io_writeReq_1_bits_data; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_1_1) begin // @[Reg.scala 17:18]
      line_write_buffer_wline_1_1 <= io_writeReq_1_bits_wline; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_1_1) begin // @[Reg.scala 17:18]
      line_write_buffer_mask_1_1 <= io_writeReq_1_bits_mask; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_1_1) begin // @[Reg.scala 17:18]
      line_write_buffer_offset_1_1 <= io_writeReq_1_bits_vwordOffset[1:0]; // @[Reg.scala 17:22]
    end
    sbuffer_in_s2_line_wen_2_1 <= io_writeReq_1_valid & io_writeReq_1_bits_wvec[2]; // @[Sbuffer.scala 131:46]
    if (sbuffer_in_s1_line_wen_2_1) begin // @[Reg.scala 17:18]
      line_write_buffer_data_2_1 <= io_writeReq_1_bits_data; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_2_1) begin // @[Reg.scala 17:18]
      line_write_buffer_wline_2_1 <= io_writeReq_1_bits_wline; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_2_1) begin // @[Reg.scala 17:18]
      line_write_buffer_mask_2_1 <= io_writeReq_1_bits_mask; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_2_1) begin // @[Reg.scala 17:18]
      line_write_buffer_offset_2_1 <= io_writeReq_1_bits_vwordOffset[1:0]; // @[Reg.scala 17:22]
    end
    sbuffer_in_s2_line_wen_3_1 <= io_writeReq_1_valid & io_writeReq_1_bits_wvec[3]; // @[Sbuffer.scala 131:46]
    if (sbuffer_in_s1_line_wen_3_1) begin // @[Reg.scala 17:18]
      line_write_buffer_data_3_1 <= io_writeReq_1_bits_data; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_3_1) begin // @[Reg.scala 17:18]
      line_write_buffer_wline_3_1 <= io_writeReq_1_bits_wline; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_3_1) begin // @[Reg.scala 17:18]
      line_write_buffer_mask_3_1 <= io_writeReq_1_bits_mask; // @[Reg.scala 17:22]
    end
    if (sbuffer_in_s1_line_wen_3_1) begin // @[Reg.scala 17:18]
      line_write_buffer_offset_3_1 <= io_writeReq_1_bits_vwordOffset[1:0]; // @[Reg.scala 17:22]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_0 <= write_byte_256 | (write_byte | _GEN_0);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_1 <= write_byte_257 | (write_byte_1 | _GEN_1);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_2 <= write_byte_258 | (write_byte_2 | _GEN_2);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_3 <= write_byte_259 | (write_byte_3 | _GEN_3);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_4 <= write_byte_260 | (write_byte_4 | _GEN_4);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_5 <= write_byte_261 | (write_byte_5 | _GEN_5);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_6 <= write_byte_262 | (write_byte_6 | _GEN_6);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_7 <= write_byte_263 | (write_byte_7 | _GEN_7);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_8 <= write_byte_264 | (write_byte_8 | _GEN_8);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_9 <= write_byte_265 | (write_byte_9 | _GEN_9);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_10 <= write_byte_266 | (write_byte_10 | _GEN_10);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_11 <= write_byte_267 | (write_byte_11 | _GEN_11);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_12 <= write_byte_268 | (write_byte_12 | _GEN_12);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_13 <= write_byte_269 | (write_byte_13 | _GEN_13);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_14 <= write_byte_270 | (write_byte_14 | _GEN_14);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_0_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_0_15 <= write_byte_271 | (write_byte_15 | _GEN_15);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_0 <= write_byte_272 | (write_byte_16 | _GEN_16);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_1 <= write_byte_273 | (write_byte_17 | _GEN_17);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_2 <= write_byte_274 | (write_byte_18 | _GEN_18);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_3 <= write_byte_275 | (write_byte_19 | _GEN_19);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_4 <= write_byte_276 | (write_byte_20 | _GEN_20);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_5 <= write_byte_277 | (write_byte_21 | _GEN_21);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_6 <= write_byte_278 | (write_byte_22 | _GEN_22);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_7 <= write_byte_279 | (write_byte_23 | _GEN_23);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_8 <= write_byte_280 | (write_byte_24 | _GEN_24);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_9 <= write_byte_281 | (write_byte_25 | _GEN_25);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_10 <= write_byte_282 | (write_byte_26 | _GEN_26);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_11 <= write_byte_283 | (write_byte_27 | _GEN_27);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_12 <= write_byte_284 | (write_byte_28 | _GEN_28);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_13 <= write_byte_285 | (write_byte_29 | _GEN_29);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_14 <= write_byte_286 | (write_byte_30 | _GEN_30);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_1_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_1_15 <= write_byte_287 | (write_byte_31 | _GEN_31);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_0 <= write_byte_288 | (write_byte_32 | _GEN_32);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_1 <= write_byte_289 | (write_byte_33 | _GEN_33);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_2 <= write_byte_290 | (write_byte_34 | _GEN_34);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_3 <= write_byte_291 | (write_byte_35 | _GEN_35);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_4 <= write_byte_292 | (write_byte_36 | _GEN_36);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_5 <= write_byte_293 | (write_byte_37 | _GEN_37);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_6 <= write_byte_294 | (write_byte_38 | _GEN_38);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_7 <= write_byte_295 | (write_byte_39 | _GEN_39);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_8 <= write_byte_296 | (write_byte_40 | _GEN_40);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_9 <= write_byte_297 | (write_byte_41 | _GEN_41);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_10 <= write_byte_298 | (write_byte_42 | _GEN_42);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_11 <= write_byte_299 | (write_byte_43 | _GEN_43);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_12 <= write_byte_300 | (write_byte_44 | _GEN_44);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_13 <= write_byte_301 | (write_byte_45 | _GEN_45);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_14 <= write_byte_302 | (write_byte_46 | _GEN_46);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_2_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_2_15 <= write_byte_303 | (write_byte_47 | _GEN_47);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_0 <= write_byte_304 | (write_byte_48 | _GEN_48);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_1 <= write_byte_305 | (write_byte_49 | _GEN_49);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_2 <= write_byte_306 | (write_byte_50 | _GEN_50);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_3 <= write_byte_307 | (write_byte_51 | _GEN_51);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_4 <= write_byte_308 | (write_byte_52 | _GEN_52);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_5 <= write_byte_309 | (write_byte_53 | _GEN_53);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_6 <= write_byte_310 | (write_byte_54 | _GEN_54);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_7 <= write_byte_311 | (write_byte_55 | _GEN_55);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_8 <= write_byte_312 | (write_byte_56 | _GEN_56);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_9 <= write_byte_313 | (write_byte_57 | _GEN_57);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_10 <= write_byte_314 | (write_byte_58 | _GEN_58);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_11 <= write_byte_315 | (write_byte_59 | _GEN_59);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_12 <= write_byte_316 | (write_byte_60 | _GEN_60);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_13 <= write_byte_317 | (write_byte_61 | _GEN_61);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_14 <= write_byte_318 | (write_byte_62 | _GEN_62);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_0_3_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_0_3_15 <= write_byte_319 | (write_byte_63 | _GEN_63);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_0 <= write_byte_320 | (write_byte_64 | _GEN_64);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_1 <= write_byte_321 | (write_byte_65 | _GEN_65);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_2 <= write_byte_322 | (write_byte_66 | _GEN_66);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_3 <= write_byte_323 | (write_byte_67 | _GEN_67);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_4 <= write_byte_324 | (write_byte_68 | _GEN_68);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_5 <= write_byte_325 | (write_byte_69 | _GEN_69);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_6 <= write_byte_326 | (write_byte_70 | _GEN_70);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_7 <= write_byte_327 | (write_byte_71 | _GEN_71);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_8 <= write_byte_328 | (write_byte_72 | _GEN_72);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_9 <= write_byte_329 | (write_byte_73 | _GEN_73);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_10 <= write_byte_330 | (write_byte_74 | _GEN_74);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_11 <= write_byte_331 | (write_byte_75 | _GEN_75);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_12 <= write_byte_332 | (write_byte_76 | _GEN_76);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_13 <= write_byte_333 | (write_byte_77 | _GEN_77);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_14 <= write_byte_334 | (write_byte_78 | _GEN_78);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_0_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_0_15 <= write_byte_335 | (write_byte_79 | _GEN_79);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_0 <= write_byte_336 | (write_byte_80 | _GEN_80);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_1 <= write_byte_337 | (write_byte_81 | _GEN_81);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_2 <= write_byte_338 | (write_byte_82 | _GEN_82);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_3 <= write_byte_339 | (write_byte_83 | _GEN_83);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_4 <= write_byte_340 | (write_byte_84 | _GEN_84);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_5 <= write_byte_341 | (write_byte_85 | _GEN_85);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_6 <= write_byte_342 | (write_byte_86 | _GEN_86);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_7 <= write_byte_343 | (write_byte_87 | _GEN_87);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_8 <= write_byte_344 | (write_byte_88 | _GEN_88);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_9 <= write_byte_345 | (write_byte_89 | _GEN_89);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_10 <= write_byte_346 | (write_byte_90 | _GEN_90);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_11 <= write_byte_347 | (write_byte_91 | _GEN_91);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_12 <= write_byte_348 | (write_byte_92 | _GEN_92);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_13 <= write_byte_349 | (write_byte_93 | _GEN_93);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_14 <= write_byte_350 | (write_byte_94 | _GEN_94);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_1_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_1_15 <= write_byte_351 | (write_byte_95 | _GEN_95);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_0 <= write_byte_352 | (write_byte_96 | _GEN_96);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_1 <= write_byte_353 | (write_byte_97 | _GEN_97);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_2 <= write_byte_354 | (write_byte_98 | _GEN_98);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_3 <= write_byte_355 | (write_byte_99 | _GEN_99);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_4 <= write_byte_356 | (write_byte_100 | _GEN_100);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_5 <= write_byte_357 | (write_byte_101 | _GEN_101);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_6 <= write_byte_358 | (write_byte_102 | _GEN_102);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_7 <= write_byte_359 | (write_byte_103 | _GEN_103);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_8 <= write_byte_360 | (write_byte_104 | _GEN_104);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_9 <= write_byte_361 | (write_byte_105 | _GEN_105);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_10 <= write_byte_362 | (write_byte_106 | _GEN_106);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_11 <= write_byte_363 | (write_byte_107 | _GEN_107);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_12 <= write_byte_364 | (write_byte_108 | _GEN_108);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_13 <= write_byte_365 | (write_byte_109 | _GEN_109);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_14 <= write_byte_366 | (write_byte_110 | _GEN_110);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_2_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_2_15 <= write_byte_367 | (write_byte_111 | _GEN_111);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_0 <= write_byte_368 | (write_byte_112 | _GEN_112);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_1 <= write_byte_369 | (write_byte_113 | _GEN_113);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_2 <= write_byte_370 | (write_byte_114 | _GEN_114);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_3 <= write_byte_371 | (write_byte_115 | _GEN_115);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_4 <= write_byte_372 | (write_byte_116 | _GEN_116);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_5 <= write_byte_373 | (write_byte_117 | _GEN_117);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_6 <= write_byte_374 | (write_byte_118 | _GEN_118);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_7 <= write_byte_375 | (write_byte_119 | _GEN_119);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_8 <= write_byte_376 | (write_byte_120 | _GEN_120);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_9 <= write_byte_377 | (write_byte_121 | _GEN_121);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_10 <= write_byte_378 | (write_byte_122 | _GEN_122);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_11 <= write_byte_379 | (write_byte_123 | _GEN_123);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_12 <= write_byte_380 | (write_byte_124 | _GEN_124);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_13 <= write_byte_381 | (write_byte_125 | _GEN_125);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_14 <= write_byte_382 | (write_byte_126 | _GEN_126);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_1_3_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_1_3_15 <= write_byte_383 | (write_byte_127 | _GEN_127);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_0 <= write_byte_384 | (write_byte_128 | _GEN_128);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_1 <= write_byte_385 | (write_byte_129 | _GEN_129);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_2 <= write_byte_386 | (write_byte_130 | _GEN_130);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_3 <= write_byte_387 | (write_byte_131 | _GEN_131);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_4 <= write_byte_388 | (write_byte_132 | _GEN_132);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_5 <= write_byte_389 | (write_byte_133 | _GEN_133);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_6 <= write_byte_390 | (write_byte_134 | _GEN_134);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_7 <= write_byte_391 | (write_byte_135 | _GEN_135);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_8 <= write_byte_392 | (write_byte_136 | _GEN_136);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_9 <= write_byte_393 | (write_byte_137 | _GEN_137);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_10 <= write_byte_394 | (write_byte_138 | _GEN_138);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_11 <= write_byte_395 | (write_byte_139 | _GEN_139);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_12 <= write_byte_396 | (write_byte_140 | _GEN_140);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_13 <= write_byte_397 | (write_byte_141 | _GEN_141);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_14 <= write_byte_398 | (write_byte_142 | _GEN_142);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_0_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_0_15 <= write_byte_399 | (write_byte_143 | _GEN_143);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_0 <= write_byte_400 | (write_byte_144 | _GEN_144);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_1 <= write_byte_401 | (write_byte_145 | _GEN_145);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_2 <= write_byte_402 | (write_byte_146 | _GEN_146);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_3 <= write_byte_403 | (write_byte_147 | _GEN_147);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_4 <= write_byte_404 | (write_byte_148 | _GEN_148);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_5 <= write_byte_405 | (write_byte_149 | _GEN_149);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_6 <= write_byte_406 | (write_byte_150 | _GEN_150);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_7 <= write_byte_407 | (write_byte_151 | _GEN_151);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_8 <= write_byte_408 | (write_byte_152 | _GEN_152);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_9 <= write_byte_409 | (write_byte_153 | _GEN_153);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_10 <= write_byte_410 | (write_byte_154 | _GEN_154);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_11 <= write_byte_411 | (write_byte_155 | _GEN_155);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_12 <= write_byte_412 | (write_byte_156 | _GEN_156);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_13 <= write_byte_413 | (write_byte_157 | _GEN_157);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_14 <= write_byte_414 | (write_byte_158 | _GEN_158);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_1_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_1_15 <= write_byte_415 | (write_byte_159 | _GEN_159);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_0 <= write_byte_416 | (write_byte_160 | _GEN_160);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_1 <= write_byte_417 | (write_byte_161 | _GEN_161);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_2 <= write_byte_418 | (write_byte_162 | _GEN_162);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_3 <= write_byte_419 | (write_byte_163 | _GEN_163);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_4 <= write_byte_420 | (write_byte_164 | _GEN_164);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_5 <= write_byte_421 | (write_byte_165 | _GEN_165);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_6 <= write_byte_422 | (write_byte_166 | _GEN_166);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_7 <= write_byte_423 | (write_byte_167 | _GEN_167);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_8 <= write_byte_424 | (write_byte_168 | _GEN_168);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_9 <= write_byte_425 | (write_byte_169 | _GEN_169);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_10 <= write_byte_426 | (write_byte_170 | _GEN_170);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_11 <= write_byte_427 | (write_byte_171 | _GEN_171);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_12 <= write_byte_428 | (write_byte_172 | _GEN_172);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_13 <= write_byte_429 | (write_byte_173 | _GEN_173);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_14 <= write_byte_430 | (write_byte_174 | _GEN_174);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_2_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_2_15 <= write_byte_431 | (write_byte_175 | _GEN_175);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_0 <= write_byte_432 | (write_byte_176 | _GEN_176);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_1 <= write_byte_433 | (write_byte_177 | _GEN_177);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_2 <= write_byte_434 | (write_byte_178 | _GEN_178);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_3 <= write_byte_435 | (write_byte_179 | _GEN_179);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_4 <= write_byte_436 | (write_byte_180 | _GEN_180);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_5 <= write_byte_437 | (write_byte_181 | _GEN_181);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_6 <= write_byte_438 | (write_byte_182 | _GEN_182);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_7 <= write_byte_439 | (write_byte_183 | _GEN_183);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_8 <= write_byte_440 | (write_byte_184 | _GEN_184);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_9 <= write_byte_441 | (write_byte_185 | _GEN_185);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_10 <= write_byte_442 | (write_byte_186 | _GEN_186);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_11 <= write_byte_443 | (write_byte_187 | _GEN_187);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_12 <= write_byte_444 | (write_byte_188 | _GEN_188);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_13 <= write_byte_445 | (write_byte_189 | _GEN_189);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_14 <= write_byte_446 | (write_byte_190 | _GEN_190);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_2_3_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_2_3_15 <= write_byte_447 | (write_byte_191 | _GEN_191);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_0 <= write_byte_448 | (write_byte_192 | _GEN_192);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_1 <= write_byte_449 | (write_byte_193 | _GEN_193);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_2 <= write_byte_450 | (write_byte_194 | _GEN_194);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_3 <= write_byte_451 | (write_byte_195 | _GEN_195);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_4 <= write_byte_452 | (write_byte_196 | _GEN_196);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_5 <= write_byte_453 | (write_byte_197 | _GEN_197);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_6 <= write_byte_454 | (write_byte_198 | _GEN_198);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_7 <= write_byte_455 | (write_byte_199 | _GEN_199);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_8 <= write_byte_456 | (write_byte_200 | _GEN_200);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_9 <= write_byte_457 | (write_byte_201 | _GEN_201);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_10 <= write_byte_458 | (write_byte_202 | _GEN_202);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_11 <= write_byte_459 | (write_byte_203 | _GEN_203);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_12 <= write_byte_460 | (write_byte_204 | _GEN_204);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_13 <= write_byte_461 | (write_byte_205 | _GEN_205);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_14 <= write_byte_462 | (write_byte_206 | _GEN_206);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_0_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_0_15 <= write_byte_463 | (write_byte_207 | _GEN_207);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_0 <= write_byte_464 | (write_byte_208 | _GEN_208);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_1 <= write_byte_465 | (write_byte_209 | _GEN_209);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_2 <= write_byte_466 | (write_byte_210 | _GEN_210);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_3 <= write_byte_467 | (write_byte_211 | _GEN_211);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_4 <= write_byte_468 | (write_byte_212 | _GEN_212);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_5 <= write_byte_469 | (write_byte_213 | _GEN_213);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_6 <= write_byte_470 | (write_byte_214 | _GEN_214);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_7 <= write_byte_471 | (write_byte_215 | _GEN_215);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_8 <= write_byte_472 | (write_byte_216 | _GEN_216);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_9 <= write_byte_473 | (write_byte_217 | _GEN_217);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_10 <= write_byte_474 | (write_byte_218 | _GEN_218);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_11 <= write_byte_475 | (write_byte_219 | _GEN_219);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_12 <= write_byte_476 | (write_byte_220 | _GEN_220);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_13 <= write_byte_477 | (write_byte_221 | _GEN_221);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_14 <= write_byte_478 | (write_byte_222 | _GEN_222);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_1_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_1_15 <= write_byte_479 | (write_byte_223 | _GEN_223);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_0 <= write_byte_480 | (write_byte_224 | _GEN_224);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_1 <= write_byte_481 | (write_byte_225 | _GEN_225);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_2 <= write_byte_482 | (write_byte_226 | _GEN_226);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_3 <= write_byte_483 | (write_byte_227 | _GEN_227);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_4 <= write_byte_484 | (write_byte_228 | _GEN_228);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_5 <= write_byte_485 | (write_byte_229 | _GEN_229);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_6 <= write_byte_486 | (write_byte_230 | _GEN_230);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_7 <= write_byte_487 | (write_byte_231 | _GEN_231);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_8 <= write_byte_488 | (write_byte_232 | _GEN_232);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_9 <= write_byte_489 | (write_byte_233 | _GEN_233);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_10 <= write_byte_490 | (write_byte_234 | _GEN_234);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_11 <= write_byte_491 | (write_byte_235 | _GEN_235);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_12 <= write_byte_492 | (write_byte_236 | _GEN_236);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_13 <= write_byte_493 | (write_byte_237 | _GEN_237);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_14 <= write_byte_494 | (write_byte_238 | _GEN_238);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_2_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_2_15 <= write_byte_495 | (write_byte_239 | _GEN_239);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_0 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_0 <= write_byte_496 | (write_byte_240 | _GEN_240);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_1 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_1 <= write_byte_497 | (write_byte_241 | _GEN_241);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_2 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_2 <= write_byte_498 | (write_byte_242 | _GEN_242);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_3 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_3 <= write_byte_499 | (write_byte_243 | _GEN_243);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_4 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_4 <= write_byte_500 | (write_byte_244 | _GEN_244);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_5 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_5 <= write_byte_501 | (write_byte_245 | _GEN_245);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_6 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_6 <= write_byte_502 | (write_byte_246 | _GEN_246);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_7 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_7 <= write_byte_503 | (write_byte_247 | _GEN_247);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_8 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_8 <= write_byte_504 | (write_byte_248 | _GEN_248);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_9 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_9 <= write_byte_505 | (write_byte_249 | _GEN_249);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_10 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_10 <= write_byte_506 | (write_byte_250 | _GEN_250);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_11 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_11 <= write_byte_507 | (write_byte_251 | _GEN_251);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_12 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_12 <= write_byte_508 | (write_byte_252 | _GEN_252);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_13 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_13 <= write_byte_509 | (write_byte_253 | _GEN_253);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_14 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_14 <= write_byte_510 | (write_byte_254 | _GEN_254);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Sbuffer.scala 149:27]
      mask_3_3_15 <= 1'h0; // @[Sbuffer.scala 151:36]
    end else begin
      mask_3_3_15 <= write_byte_511 | (write_byte_255 | _GEN_255);
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_0_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_0_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_0_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_0_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_0_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_0_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_0_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_0_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_0_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_0_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_0_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_0_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_1_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_1_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_1_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_1_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_1_4 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_1_5 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_1_6 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_1_7 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_1_8 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_1_9 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_1_10 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_1_11 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_1_12 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_1_13 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_1_14 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_1_15 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_0_2_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_0_2_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_0_2_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_0_2_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_0_2_4 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_0_2_5 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_0_2_6 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_0_2_7 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_0_2_8 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_0_2_9 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_0_2_10 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_0_2_11 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_0_2_12 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_0_2_13 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_0_2_14 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_0_2_15 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_0_3_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_0_3_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_0_3_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_0_3_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_0_3_4 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_0_3_5 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_0_3_6 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_0_3_7 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_0_3_8 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_0_3_9 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_0_3_10 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_0_3_11 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_0_3_12 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_0_3_13 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_0_3_14 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_0_3_15 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  data_1_0_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  data_1_0_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  data_1_0_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  data_1_0_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  data_1_0_4 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  data_1_0_5 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  data_1_0_6 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  data_1_0_7 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  data_1_0_8 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  data_1_0_9 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  data_1_0_10 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  data_1_0_11 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  data_1_0_12 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  data_1_0_13 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  data_1_0_14 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  data_1_0_15 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  data_1_1_0 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  data_1_1_1 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  data_1_1_2 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  data_1_1_3 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  data_1_1_4 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  data_1_1_5 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  data_1_1_6 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  data_1_1_7 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  data_1_1_8 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  data_1_1_9 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  data_1_1_10 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  data_1_1_11 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  data_1_1_12 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  data_1_1_13 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  data_1_1_14 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  data_1_1_15 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  data_1_2_0 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  data_1_2_1 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  data_1_2_2 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  data_1_2_3 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  data_1_2_4 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  data_1_2_5 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  data_1_2_6 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  data_1_2_7 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  data_1_2_8 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  data_1_2_9 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  data_1_2_10 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  data_1_2_11 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  data_1_2_12 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  data_1_2_13 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  data_1_2_14 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  data_1_2_15 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  data_1_3_0 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  data_1_3_1 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  data_1_3_2 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  data_1_3_3 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  data_1_3_4 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  data_1_3_5 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  data_1_3_6 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  data_1_3_7 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  data_1_3_8 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  data_1_3_9 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  data_1_3_10 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  data_1_3_11 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  data_1_3_12 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  data_1_3_13 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  data_1_3_14 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  data_1_3_15 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  data_2_0_0 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  data_2_0_1 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  data_2_0_2 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  data_2_0_3 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  data_2_0_4 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  data_2_0_5 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  data_2_0_6 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  data_2_0_7 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  data_2_0_8 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  data_2_0_9 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  data_2_0_10 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  data_2_0_11 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  data_2_0_12 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  data_2_0_13 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  data_2_0_14 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  data_2_0_15 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  data_2_1_0 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  data_2_1_1 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  data_2_1_2 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  data_2_1_3 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  data_2_1_4 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  data_2_1_5 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  data_2_1_6 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  data_2_1_7 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  data_2_1_8 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  data_2_1_9 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  data_2_1_10 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  data_2_1_11 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  data_2_1_12 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  data_2_1_13 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  data_2_1_14 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  data_2_1_15 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  data_2_2_0 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  data_2_2_1 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  data_2_2_2 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  data_2_2_3 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  data_2_2_4 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  data_2_2_5 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  data_2_2_6 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  data_2_2_7 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  data_2_2_8 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  data_2_2_9 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  data_2_2_10 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  data_2_2_11 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  data_2_2_12 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  data_2_2_13 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  data_2_2_14 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  data_2_2_15 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  data_2_3_0 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  data_2_3_1 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  data_2_3_2 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  data_2_3_3 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  data_2_3_4 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  data_2_3_5 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  data_2_3_6 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  data_2_3_7 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  data_2_3_8 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  data_2_3_9 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  data_2_3_10 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  data_2_3_11 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  data_2_3_12 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  data_2_3_13 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  data_2_3_14 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  data_2_3_15 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  data_3_0_0 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  data_3_0_1 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  data_3_0_2 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  data_3_0_3 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  data_3_0_4 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  data_3_0_5 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  data_3_0_6 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  data_3_0_7 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  data_3_0_8 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  data_3_0_9 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  data_3_0_10 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  data_3_0_11 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  data_3_0_12 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  data_3_0_13 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  data_3_0_14 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  data_3_0_15 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  data_3_1_0 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  data_3_1_1 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  data_3_1_2 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  data_3_1_3 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  data_3_1_4 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  data_3_1_5 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  data_3_1_6 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  data_3_1_7 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  data_3_1_8 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  data_3_1_9 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  data_3_1_10 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  data_3_1_11 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  data_3_1_12 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  data_3_1_13 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  data_3_1_14 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  data_3_1_15 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  data_3_2_0 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  data_3_2_1 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  data_3_2_2 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  data_3_2_3 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  data_3_2_4 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  data_3_2_5 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  data_3_2_6 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  data_3_2_7 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  data_3_2_8 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  data_3_2_9 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  data_3_2_10 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  data_3_2_11 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  data_3_2_12 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  data_3_2_13 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  data_3_2_14 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  data_3_2_15 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  data_3_3_0 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  data_3_3_1 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  data_3_3_2 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  data_3_3_3 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  data_3_3_4 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  data_3_3_5 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  data_3_3_6 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  data_3_3_7 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  data_3_3_8 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  data_3_3_9 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  data_3_3_10 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  data_3_3_11 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  data_3_3_12 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  data_3_3_13 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  data_3_3_14 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  data_3_3_15 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  mask_0_0_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  mask_0_0_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  mask_0_0_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  mask_0_0_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  mask_0_0_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  mask_0_0_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  mask_0_0_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  mask_0_0_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  mask_0_0_8 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  mask_0_0_9 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  mask_0_0_10 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  mask_0_0_11 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  mask_0_0_12 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  mask_0_0_13 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  mask_0_0_14 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  mask_0_0_15 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  mask_0_1_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  mask_0_1_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  mask_0_1_2 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  mask_0_1_3 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  mask_0_1_4 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  mask_0_1_5 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  mask_0_1_6 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  mask_0_1_7 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  mask_0_1_8 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  mask_0_1_9 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  mask_0_1_10 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  mask_0_1_11 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  mask_0_1_12 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  mask_0_1_13 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  mask_0_1_14 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  mask_0_1_15 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  mask_0_2_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  mask_0_2_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  mask_0_2_2 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  mask_0_2_3 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  mask_0_2_4 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  mask_0_2_5 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  mask_0_2_6 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  mask_0_2_7 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  mask_0_2_8 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  mask_0_2_9 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  mask_0_2_10 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  mask_0_2_11 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  mask_0_2_12 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  mask_0_2_13 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  mask_0_2_14 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  mask_0_2_15 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  mask_0_3_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  mask_0_3_1 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  mask_0_3_2 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  mask_0_3_3 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  mask_0_3_4 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  mask_0_3_5 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  mask_0_3_6 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  mask_0_3_7 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  mask_0_3_8 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  mask_0_3_9 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  mask_0_3_10 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  mask_0_3_11 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  mask_0_3_12 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  mask_0_3_13 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  mask_0_3_14 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  mask_0_3_15 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  mask_1_0_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  mask_1_0_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  mask_1_0_2 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  mask_1_0_3 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  mask_1_0_4 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  mask_1_0_5 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  mask_1_0_6 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  mask_1_0_7 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  mask_1_0_8 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  mask_1_0_9 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  mask_1_0_10 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  mask_1_0_11 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  mask_1_0_12 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  mask_1_0_13 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  mask_1_0_14 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  mask_1_0_15 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  mask_1_1_0 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  mask_1_1_1 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  mask_1_1_2 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  mask_1_1_3 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  mask_1_1_4 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  mask_1_1_5 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  mask_1_1_6 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  mask_1_1_7 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  mask_1_1_8 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  mask_1_1_9 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  mask_1_1_10 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  mask_1_1_11 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  mask_1_1_12 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  mask_1_1_13 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  mask_1_1_14 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  mask_1_1_15 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  mask_1_2_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  mask_1_2_1 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  mask_1_2_2 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  mask_1_2_3 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  mask_1_2_4 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  mask_1_2_5 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  mask_1_2_6 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  mask_1_2_7 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  mask_1_2_8 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  mask_1_2_9 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  mask_1_2_10 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  mask_1_2_11 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  mask_1_2_12 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  mask_1_2_13 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  mask_1_2_14 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  mask_1_2_15 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  mask_1_3_0 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  mask_1_3_1 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  mask_1_3_2 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  mask_1_3_3 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  mask_1_3_4 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  mask_1_3_5 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  mask_1_3_6 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  mask_1_3_7 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  mask_1_3_8 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  mask_1_3_9 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  mask_1_3_10 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  mask_1_3_11 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  mask_1_3_12 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  mask_1_3_13 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  mask_1_3_14 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  mask_1_3_15 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  mask_2_0_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  mask_2_0_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  mask_2_0_2 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  mask_2_0_3 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  mask_2_0_4 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  mask_2_0_5 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  mask_2_0_6 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  mask_2_0_7 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  mask_2_0_8 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  mask_2_0_9 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  mask_2_0_10 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  mask_2_0_11 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  mask_2_0_12 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  mask_2_0_13 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  mask_2_0_14 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  mask_2_0_15 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  mask_2_1_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  mask_2_1_1 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  mask_2_1_2 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  mask_2_1_3 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  mask_2_1_4 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  mask_2_1_5 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  mask_2_1_6 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  mask_2_1_7 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  mask_2_1_8 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  mask_2_1_9 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  mask_2_1_10 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  mask_2_1_11 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  mask_2_1_12 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  mask_2_1_13 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  mask_2_1_14 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  mask_2_1_15 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  mask_2_2_0 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  mask_2_2_1 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  mask_2_2_2 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  mask_2_2_3 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  mask_2_2_4 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  mask_2_2_5 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  mask_2_2_6 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  mask_2_2_7 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  mask_2_2_8 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  mask_2_2_9 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  mask_2_2_10 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  mask_2_2_11 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  mask_2_2_12 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  mask_2_2_13 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  mask_2_2_14 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  mask_2_2_15 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  mask_2_3_0 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  mask_2_3_1 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  mask_2_3_2 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  mask_2_3_3 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  mask_2_3_4 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  mask_2_3_5 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  mask_2_3_6 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  mask_2_3_7 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  mask_2_3_8 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  mask_2_3_9 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  mask_2_3_10 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  mask_2_3_11 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  mask_2_3_12 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  mask_2_3_13 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  mask_2_3_14 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  mask_2_3_15 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  mask_3_0_0 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  mask_3_0_1 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  mask_3_0_2 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  mask_3_0_3 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  mask_3_0_4 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  mask_3_0_5 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  mask_3_0_6 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  mask_3_0_7 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  mask_3_0_8 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  mask_3_0_9 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  mask_3_0_10 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  mask_3_0_11 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  mask_3_0_12 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  mask_3_0_13 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  mask_3_0_14 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  mask_3_0_15 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  mask_3_1_0 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  mask_3_1_1 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  mask_3_1_2 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  mask_3_1_3 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  mask_3_1_4 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  mask_3_1_5 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  mask_3_1_6 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  mask_3_1_7 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  mask_3_1_8 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  mask_3_1_9 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  mask_3_1_10 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  mask_3_1_11 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  mask_3_1_12 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  mask_3_1_13 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  mask_3_1_14 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  mask_3_1_15 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  mask_3_2_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  mask_3_2_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  mask_3_2_2 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  mask_3_2_3 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  mask_3_2_4 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  mask_3_2_5 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  mask_3_2_6 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  mask_3_2_7 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  mask_3_2_8 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  mask_3_2_9 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  mask_3_2_10 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  mask_3_2_11 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  mask_3_2_12 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  mask_3_2_13 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  mask_3_2_14 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  mask_3_2_15 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  mask_3_3_0 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  mask_3_3_1 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  mask_3_3_2 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  mask_3_3_3 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  mask_3_3_4 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  mask_3_3_5 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  mask_3_3_6 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  mask_3_3_7 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  mask_3_3_8 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  mask_3_3_9 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  mask_3_3_10 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  mask_3_3_11 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  mask_3_3_12 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  mask_3_3_13 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  mask_3_3_14 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  mask_3_3_15 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  line_mask_clean_flag_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  line_mask_clean_flag_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  line_mask_clean_flag_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  line_mask_clean_flag_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  sbuffer_in_s2_line_wen_0 = _RAND_516[0:0];
  _RAND_517 = {4{`RANDOM}};
  line_write_buffer_data_0 = _RAND_517[127:0];
  _RAND_518 = {1{`RANDOM}};
  line_write_buffer_wline_0 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  line_write_buffer_mask_0 = _RAND_519[15:0];
  _RAND_520 = {1{`RANDOM}};
  line_write_buffer_offset_0 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  sbuffer_in_s2_line_wen_1 = _RAND_521[0:0];
  _RAND_522 = {4{`RANDOM}};
  line_write_buffer_data_1 = _RAND_522[127:0];
  _RAND_523 = {1{`RANDOM}};
  line_write_buffer_wline_1 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  line_write_buffer_mask_1 = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  line_write_buffer_offset_1 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  sbuffer_in_s2_line_wen_2 = _RAND_526[0:0];
  _RAND_527 = {4{`RANDOM}};
  line_write_buffer_data_2 = _RAND_527[127:0];
  _RAND_528 = {1{`RANDOM}};
  line_write_buffer_wline_2 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  line_write_buffer_mask_2 = _RAND_529[15:0];
  _RAND_530 = {1{`RANDOM}};
  line_write_buffer_offset_2 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  sbuffer_in_s2_line_wen_3 = _RAND_531[0:0];
  _RAND_532 = {4{`RANDOM}};
  line_write_buffer_data_3 = _RAND_532[127:0];
  _RAND_533 = {1{`RANDOM}};
  line_write_buffer_wline_3 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  line_write_buffer_mask_3 = _RAND_534[15:0];
  _RAND_535 = {1{`RANDOM}};
  line_write_buffer_offset_3 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  sbuffer_in_s2_line_wen_0_1 = _RAND_536[0:0];
  _RAND_537 = {4{`RANDOM}};
  line_write_buffer_data_0_1 = _RAND_537[127:0];
  _RAND_538 = {1{`RANDOM}};
  line_write_buffer_wline_0_1 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  line_write_buffer_mask_0_1 = _RAND_539[15:0];
  _RAND_540 = {1{`RANDOM}};
  line_write_buffer_offset_0_1 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  sbuffer_in_s2_line_wen_1_1 = _RAND_541[0:0];
  _RAND_542 = {4{`RANDOM}};
  line_write_buffer_data_1_1 = _RAND_542[127:0];
  _RAND_543 = {1{`RANDOM}};
  line_write_buffer_wline_1_1 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  line_write_buffer_mask_1_1 = _RAND_544[15:0];
  _RAND_545 = {1{`RANDOM}};
  line_write_buffer_offset_1_1 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  sbuffer_in_s2_line_wen_2_1 = _RAND_546[0:0];
  _RAND_547 = {4{`RANDOM}};
  line_write_buffer_data_2_1 = _RAND_547[127:0];
  _RAND_548 = {1{`RANDOM}};
  line_write_buffer_wline_2_1 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  line_write_buffer_mask_2_1 = _RAND_549[15:0];
  _RAND_550 = {1{`RANDOM}};
  line_write_buffer_offset_2_1 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  sbuffer_in_s2_line_wen_3_1 = _RAND_551[0:0];
  _RAND_552 = {4{`RANDOM}};
  line_write_buffer_data_3_1 = _RAND_552[127:0];
  _RAND_553 = {1{`RANDOM}};
  line_write_buffer_wline_3_1 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  line_write_buffer_mask_3_1 = _RAND_554[15:0];
  _RAND_555 = {1{`RANDOM}};
  line_write_buffer_offset_3_1 = _RAND_555[1:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    mask_0_0_0 = 1'h0;
  end
  if (reset) begin
    mask_0_0_1 = 1'h0;
  end
  if (reset) begin
    mask_0_0_2 = 1'h0;
  end
  if (reset) begin
    mask_0_0_3 = 1'h0;
  end
  if (reset) begin
    mask_0_0_4 = 1'h0;
  end
  if (reset) begin
    mask_0_0_5 = 1'h0;
  end
  if (reset) begin
    mask_0_0_6 = 1'h0;
  end
  if (reset) begin
    mask_0_0_7 = 1'h0;
  end
  if (reset) begin
    mask_0_0_8 = 1'h0;
  end
  if (reset) begin
    mask_0_0_9 = 1'h0;
  end
  if (reset) begin
    mask_0_0_10 = 1'h0;
  end
  if (reset) begin
    mask_0_0_11 = 1'h0;
  end
  if (reset) begin
    mask_0_0_12 = 1'h0;
  end
  if (reset) begin
    mask_0_0_13 = 1'h0;
  end
  if (reset) begin
    mask_0_0_14 = 1'h0;
  end
  if (reset) begin
    mask_0_0_15 = 1'h0;
  end
  if (reset) begin
    mask_0_1_0 = 1'h0;
  end
  if (reset) begin
    mask_0_1_1 = 1'h0;
  end
  if (reset) begin
    mask_0_1_2 = 1'h0;
  end
  if (reset) begin
    mask_0_1_3 = 1'h0;
  end
  if (reset) begin
    mask_0_1_4 = 1'h0;
  end
  if (reset) begin
    mask_0_1_5 = 1'h0;
  end
  if (reset) begin
    mask_0_1_6 = 1'h0;
  end
  if (reset) begin
    mask_0_1_7 = 1'h0;
  end
  if (reset) begin
    mask_0_1_8 = 1'h0;
  end
  if (reset) begin
    mask_0_1_9 = 1'h0;
  end
  if (reset) begin
    mask_0_1_10 = 1'h0;
  end
  if (reset) begin
    mask_0_1_11 = 1'h0;
  end
  if (reset) begin
    mask_0_1_12 = 1'h0;
  end
  if (reset) begin
    mask_0_1_13 = 1'h0;
  end
  if (reset) begin
    mask_0_1_14 = 1'h0;
  end
  if (reset) begin
    mask_0_1_15 = 1'h0;
  end
  if (reset) begin
    mask_0_2_0 = 1'h0;
  end
  if (reset) begin
    mask_0_2_1 = 1'h0;
  end
  if (reset) begin
    mask_0_2_2 = 1'h0;
  end
  if (reset) begin
    mask_0_2_3 = 1'h0;
  end
  if (reset) begin
    mask_0_2_4 = 1'h0;
  end
  if (reset) begin
    mask_0_2_5 = 1'h0;
  end
  if (reset) begin
    mask_0_2_6 = 1'h0;
  end
  if (reset) begin
    mask_0_2_7 = 1'h0;
  end
  if (reset) begin
    mask_0_2_8 = 1'h0;
  end
  if (reset) begin
    mask_0_2_9 = 1'h0;
  end
  if (reset) begin
    mask_0_2_10 = 1'h0;
  end
  if (reset) begin
    mask_0_2_11 = 1'h0;
  end
  if (reset) begin
    mask_0_2_12 = 1'h0;
  end
  if (reset) begin
    mask_0_2_13 = 1'h0;
  end
  if (reset) begin
    mask_0_2_14 = 1'h0;
  end
  if (reset) begin
    mask_0_2_15 = 1'h0;
  end
  if (reset) begin
    mask_0_3_0 = 1'h0;
  end
  if (reset) begin
    mask_0_3_1 = 1'h0;
  end
  if (reset) begin
    mask_0_3_2 = 1'h0;
  end
  if (reset) begin
    mask_0_3_3 = 1'h0;
  end
  if (reset) begin
    mask_0_3_4 = 1'h0;
  end
  if (reset) begin
    mask_0_3_5 = 1'h0;
  end
  if (reset) begin
    mask_0_3_6 = 1'h0;
  end
  if (reset) begin
    mask_0_3_7 = 1'h0;
  end
  if (reset) begin
    mask_0_3_8 = 1'h0;
  end
  if (reset) begin
    mask_0_3_9 = 1'h0;
  end
  if (reset) begin
    mask_0_3_10 = 1'h0;
  end
  if (reset) begin
    mask_0_3_11 = 1'h0;
  end
  if (reset) begin
    mask_0_3_12 = 1'h0;
  end
  if (reset) begin
    mask_0_3_13 = 1'h0;
  end
  if (reset) begin
    mask_0_3_14 = 1'h0;
  end
  if (reset) begin
    mask_0_3_15 = 1'h0;
  end
  if (reset) begin
    mask_1_0_0 = 1'h0;
  end
  if (reset) begin
    mask_1_0_1 = 1'h0;
  end
  if (reset) begin
    mask_1_0_2 = 1'h0;
  end
  if (reset) begin
    mask_1_0_3 = 1'h0;
  end
  if (reset) begin
    mask_1_0_4 = 1'h0;
  end
  if (reset) begin
    mask_1_0_5 = 1'h0;
  end
  if (reset) begin
    mask_1_0_6 = 1'h0;
  end
  if (reset) begin
    mask_1_0_7 = 1'h0;
  end
  if (reset) begin
    mask_1_0_8 = 1'h0;
  end
  if (reset) begin
    mask_1_0_9 = 1'h0;
  end
  if (reset) begin
    mask_1_0_10 = 1'h0;
  end
  if (reset) begin
    mask_1_0_11 = 1'h0;
  end
  if (reset) begin
    mask_1_0_12 = 1'h0;
  end
  if (reset) begin
    mask_1_0_13 = 1'h0;
  end
  if (reset) begin
    mask_1_0_14 = 1'h0;
  end
  if (reset) begin
    mask_1_0_15 = 1'h0;
  end
  if (reset) begin
    mask_1_1_0 = 1'h0;
  end
  if (reset) begin
    mask_1_1_1 = 1'h0;
  end
  if (reset) begin
    mask_1_1_2 = 1'h0;
  end
  if (reset) begin
    mask_1_1_3 = 1'h0;
  end
  if (reset) begin
    mask_1_1_4 = 1'h0;
  end
  if (reset) begin
    mask_1_1_5 = 1'h0;
  end
  if (reset) begin
    mask_1_1_6 = 1'h0;
  end
  if (reset) begin
    mask_1_1_7 = 1'h0;
  end
  if (reset) begin
    mask_1_1_8 = 1'h0;
  end
  if (reset) begin
    mask_1_1_9 = 1'h0;
  end
  if (reset) begin
    mask_1_1_10 = 1'h0;
  end
  if (reset) begin
    mask_1_1_11 = 1'h0;
  end
  if (reset) begin
    mask_1_1_12 = 1'h0;
  end
  if (reset) begin
    mask_1_1_13 = 1'h0;
  end
  if (reset) begin
    mask_1_1_14 = 1'h0;
  end
  if (reset) begin
    mask_1_1_15 = 1'h0;
  end
  if (reset) begin
    mask_1_2_0 = 1'h0;
  end
  if (reset) begin
    mask_1_2_1 = 1'h0;
  end
  if (reset) begin
    mask_1_2_2 = 1'h0;
  end
  if (reset) begin
    mask_1_2_3 = 1'h0;
  end
  if (reset) begin
    mask_1_2_4 = 1'h0;
  end
  if (reset) begin
    mask_1_2_5 = 1'h0;
  end
  if (reset) begin
    mask_1_2_6 = 1'h0;
  end
  if (reset) begin
    mask_1_2_7 = 1'h0;
  end
  if (reset) begin
    mask_1_2_8 = 1'h0;
  end
  if (reset) begin
    mask_1_2_9 = 1'h0;
  end
  if (reset) begin
    mask_1_2_10 = 1'h0;
  end
  if (reset) begin
    mask_1_2_11 = 1'h0;
  end
  if (reset) begin
    mask_1_2_12 = 1'h0;
  end
  if (reset) begin
    mask_1_2_13 = 1'h0;
  end
  if (reset) begin
    mask_1_2_14 = 1'h0;
  end
  if (reset) begin
    mask_1_2_15 = 1'h0;
  end
  if (reset) begin
    mask_1_3_0 = 1'h0;
  end
  if (reset) begin
    mask_1_3_1 = 1'h0;
  end
  if (reset) begin
    mask_1_3_2 = 1'h0;
  end
  if (reset) begin
    mask_1_3_3 = 1'h0;
  end
  if (reset) begin
    mask_1_3_4 = 1'h0;
  end
  if (reset) begin
    mask_1_3_5 = 1'h0;
  end
  if (reset) begin
    mask_1_3_6 = 1'h0;
  end
  if (reset) begin
    mask_1_3_7 = 1'h0;
  end
  if (reset) begin
    mask_1_3_8 = 1'h0;
  end
  if (reset) begin
    mask_1_3_9 = 1'h0;
  end
  if (reset) begin
    mask_1_3_10 = 1'h0;
  end
  if (reset) begin
    mask_1_3_11 = 1'h0;
  end
  if (reset) begin
    mask_1_3_12 = 1'h0;
  end
  if (reset) begin
    mask_1_3_13 = 1'h0;
  end
  if (reset) begin
    mask_1_3_14 = 1'h0;
  end
  if (reset) begin
    mask_1_3_15 = 1'h0;
  end
  if (reset) begin
    mask_2_0_0 = 1'h0;
  end
  if (reset) begin
    mask_2_0_1 = 1'h0;
  end
  if (reset) begin
    mask_2_0_2 = 1'h0;
  end
  if (reset) begin
    mask_2_0_3 = 1'h0;
  end
  if (reset) begin
    mask_2_0_4 = 1'h0;
  end
  if (reset) begin
    mask_2_0_5 = 1'h0;
  end
  if (reset) begin
    mask_2_0_6 = 1'h0;
  end
  if (reset) begin
    mask_2_0_7 = 1'h0;
  end
  if (reset) begin
    mask_2_0_8 = 1'h0;
  end
  if (reset) begin
    mask_2_0_9 = 1'h0;
  end
  if (reset) begin
    mask_2_0_10 = 1'h0;
  end
  if (reset) begin
    mask_2_0_11 = 1'h0;
  end
  if (reset) begin
    mask_2_0_12 = 1'h0;
  end
  if (reset) begin
    mask_2_0_13 = 1'h0;
  end
  if (reset) begin
    mask_2_0_14 = 1'h0;
  end
  if (reset) begin
    mask_2_0_15 = 1'h0;
  end
  if (reset) begin
    mask_2_1_0 = 1'h0;
  end
  if (reset) begin
    mask_2_1_1 = 1'h0;
  end
  if (reset) begin
    mask_2_1_2 = 1'h0;
  end
  if (reset) begin
    mask_2_1_3 = 1'h0;
  end
  if (reset) begin
    mask_2_1_4 = 1'h0;
  end
  if (reset) begin
    mask_2_1_5 = 1'h0;
  end
  if (reset) begin
    mask_2_1_6 = 1'h0;
  end
  if (reset) begin
    mask_2_1_7 = 1'h0;
  end
  if (reset) begin
    mask_2_1_8 = 1'h0;
  end
  if (reset) begin
    mask_2_1_9 = 1'h0;
  end
  if (reset) begin
    mask_2_1_10 = 1'h0;
  end
  if (reset) begin
    mask_2_1_11 = 1'h0;
  end
  if (reset) begin
    mask_2_1_12 = 1'h0;
  end
  if (reset) begin
    mask_2_1_13 = 1'h0;
  end
  if (reset) begin
    mask_2_1_14 = 1'h0;
  end
  if (reset) begin
    mask_2_1_15 = 1'h0;
  end
  if (reset) begin
    mask_2_2_0 = 1'h0;
  end
  if (reset) begin
    mask_2_2_1 = 1'h0;
  end
  if (reset) begin
    mask_2_2_2 = 1'h0;
  end
  if (reset) begin
    mask_2_2_3 = 1'h0;
  end
  if (reset) begin
    mask_2_2_4 = 1'h0;
  end
  if (reset) begin
    mask_2_2_5 = 1'h0;
  end
  if (reset) begin
    mask_2_2_6 = 1'h0;
  end
  if (reset) begin
    mask_2_2_7 = 1'h0;
  end
  if (reset) begin
    mask_2_2_8 = 1'h0;
  end
  if (reset) begin
    mask_2_2_9 = 1'h0;
  end
  if (reset) begin
    mask_2_2_10 = 1'h0;
  end
  if (reset) begin
    mask_2_2_11 = 1'h0;
  end
  if (reset) begin
    mask_2_2_12 = 1'h0;
  end
  if (reset) begin
    mask_2_2_13 = 1'h0;
  end
  if (reset) begin
    mask_2_2_14 = 1'h0;
  end
  if (reset) begin
    mask_2_2_15 = 1'h0;
  end
  if (reset) begin
    mask_2_3_0 = 1'h0;
  end
  if (reset) begin
    mask_2_3_1 = 1'h0;
  end
  if (reset) begin
    mask_2_3_2 = 1'h0;
  end
  if (reset) begin
    mask_2_3_3 = 1'h0;
  end
  if (reset) begin
    mask_2_3_4 = 1'h0;
  end
  if (reset) begin
    mask_2_3_5 = 1'h0;
  end
  if (reset) begin
    mask_2_3_6 = 1'h0;
  end
  if (reset) begin
    mask_2_3_7 = 1'h0;
  end
  if (reset) begin
    mask_2_3_8 = 1'h0;
  end
  if (reset) begin
    mask_2_3_9 = 1'h0;
  end
  if (reset) begin
    mask_2_3_10 = 1'h0;
  end
  if (reset) begin
    mask_2_3_11 = 1'h0;
  end
  if (reset) begin
    mask_2_3_12 = 1'h0;
  end
  if (reset) begin
    mask_2_3_13 = 1'h0;
  end
  if (reset) begin
    mask_2_3_14 = 1'h0;
  end
  if (reset) begin
    mask_2_3_15 = 1'h0;
  end
  if (reset) begin
    mask_3_0_0 = 1'h0;
  end
  if (reset) begin
    mask_3_0_1 = 1'h0;
  end
  if (reset) begin
    mask_3_0_2 = 1'h0;
  end
  if (reset) begin
    mask_3_0_3 = 1'h0;
  end
  if (reset) begin
    mask_3_0_4 = 1'h0;
  end
  if (reset) begin
    mask_3_0_5 = 1'h0;
  end
  if (reset) begin
    mask_3_0_6 = 1'h0;
  end
  if (reset) begin
    mask_3_0_7 = 1'h0;
  end
  if (reset) begin
    mask_3_0_8 = 1'h0;
  end
  if (reset) begin
    mask_3_0_9 = 1'h0;
  end
  if (reset) begin
    mask_3_0_10 = 1'h0;
  end
  if (reset) begin
    mask_3_0_11 = 1'h0;
  end
  if (reset) begin
    mask_3_0_12 = 1'h0;
  end
  if (reset) begin
    mask_3_0_13 = 1'h0;
  end
  if (reset) begin
    mask_3_0_14 = 1'h0;
  end
  if (reset) begin
    mask_3_0_15 = 1'h0;
  end
  if (reset) begin
    mask_3_1_0 = 1'h0;
  end
  if (reset) begin
    mask_3_1_1 = 1'h0;
  end
  if (reset) begin
    mask_3_1_2 = 1'h0;
  end
  if (reset) begin
    mask_3_1_3 = 1'h0;
  end
  if (reset) begin
    mask_3_1_4 = 1'h0;
  end
  if (reset) begin
    mask_3_1_5 = 1'h0;
  end
  if (reset) begin
    mask_3_1_6 = 1'h0;
  end
  if (reset) begin
    mask_3_1_7 = 1'h0;
  end
  if (reset) begin
    mask_3_1_8 = 1'h0;
  end
  if (reset) begin
    mask_3_1_9 = 1'h0;
  end
  if (reset) begin
    mask_3_1_10 = 1'h0;
  end
  if (reset) begin
    mask_3_1_11 = 1'h0;
  end
  if (reset) begin
    mask_3_1_12 = 1'h0;
  end
  if (reset) begin
    mask_3_1_13 = 1'h0;
  end
  if (reset) begin
    mask_3_1_14 = 1'h0;
  end
  if (reset) begin
    mask_3_1_15 = 1'h0;
  end
  if (reset) begin
    mask_3_2_0 = 1'h0;
  end
  if (reset) begin
    mask_3_2_1 = 1'h0;
  end
  if (reset) begin
    mask_3_2_2 = 1'h0;
  end
  if (reset) begin
    mask_3_2_3 = 1'h0;
  end
  if (reset) begin
    mask_3_2_4 = 1'h0;
  end
  if (reset) begin
    mask_3_2_5 = 1'h0;
  end
  if (reset) begin
    mask_3_2_6 = 1'h0;
  end
  if (reset) begin
    mask_3_2_7 = 1'h0;
  end
  if (reset) begin
    mask_3_2_8 = 1'h0;
  end
  if (reset) begin
    mask_3_2_9 = 1'h0;
  end
  if (reset) begin
    mask_3_2_10 = 1'h0;
  end
  if (reset) begin
    mask_3_2_11 = 1'h0;
  end
  if (reset) begin
    mask_3_2_12 = 1'h0;
  end
  if (reset) begin
    mask_3_2_13 = 1'h0;
  end
  if (reset) begin
    mask_3_2_14 = 1'h0;
  end
  if (reset) begin
    mask_3_2_15 = 1'h0;
  end
  if (reset) begin
    mask_3_3_0 = 1'h0;
  end
  if (reset) begin
    mask_3_3_1 = 1'h0;
  end
  if (reset) begin
    mask_3_3_2 = 1'h0;
  end
  if (reset) begin
    mask_3_3_3 = 1'h0;
  end
  if (reset) begin
    mask_3_3_4 = 1'h0;
  end
  if (reset) begin
    mask_3_3_5 = 1'h0;
  end
  if (reset) begin
    mask_3_3_6 = 1'h0;
  end
  if (reset) begin
    mask_3_3_7 = 1'h0;
  end
  if (reset) begin
    mask_3_3_8 = 1'h0;
  end
  if (reset) begin
    mask_3_3_9 = 1'h0;
  end
  if (reset) begin
    mask_3_3_10 = 1'h0;
  end
  if (reset) begin
    mask_3_3_11 = 1'h0;
  end
  if (reset) begin
    mask_3_3_12 = 1'h0;
  end
  if (reset) begin
    mask_3_3_13 = 1'h0;
  end
  if (reset) begin
    mask_3_3_14 = 1'h0;
  end
  if (reset) begin
    mask_3_3_15 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

