module ITTageTable_3(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [38:0] io_req_bits_pc,
  input  [8:0]  io_req_bits_folded_hist_hist_7_folded_hist,
  input  [7:0]  io_req_bits_folded_hist_hist_0_folded_hist,
  output        io_resp_valid,
  output [1:0]  io_resp_bits_ctr,
  output [1:0]  io_resp_bits_u,
  output [38:0] io_resp_bits_target,
  input  [38:0] io_update_pc,
  input  [8:0]  io_update_folded_hist_hist_7_folded_hist,
  input  [7:0]  io_update_folded_hist_hist_0_folded_hist,
  input         io_update_valid,
  input         io_update_correct,
  input         io_update_alloc,
  input  [1:0]  io_update_oldCtr,
  input         io_update_uValid,
  input         io_update_u,
  input         io_update_reset_u,
  input  [38:0] io_update_target,
  input  [38:0] io_update_old_target
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  us_clock; // @[ITTAGE.scala 222:18]
  wire  us_reset; // @[ITTAGE.scala 222:18]
  wire [8:0] us_io_raddr_0; // @[ITTAGE.scala 222:18]
  wire  us_io_rdata_0; // @[ITTAGE.scala 222:18]
  wire  us_io_wen; // @[ITTAGE.scala 222:18]
  wire [8:0] us_io_waddr; // @[ITTAGE.scala 222:18]
  wire  us_io_wdata; // @[ITTAGE.scala 222:18]
  wire  us_io_resetEn; // @[ITTAGE.scala 222:18]
  wire  table_banks_0_clock; // @[ITTAGE.scala 225:11]
  wire  table_banks_0_reset; // @[ITTAGE.scala 225:11]
  wire  table_banks_0_io_rreq_valid; // @[ITTAGE.scala 225:11]
  wire [7:0] table_banks_0_io_rreq_bits_setIdx; // @[ITTAGE.scala 225:11]
  wire [8:0] table_banks_0_io_rresp_data_0_tag; // @[ITTAGE.scala 225:11]
  wire [1:0] table_banks_0_io_rresp_data_0_ctr; // @[ITTAGE.scala 225:11]
  wire [38:0] table_banks_0_io_rresp_data_0_target; // @[ITTAGE.scala 225:11]
  wire  table_banks_0_io_wreq_valid; // @[ITTAGE.scala 225:11]
  wire [7:0] table_banks_0_io_wreq_bits_setIdx; // @[ITTAGE.scala 225:11]
  wire [8:0] table_banks_0_io_wreq_bits_data_0_tag; // @[ITTAGE.scala 225:11]
  wire [1:0] table_banks_0_io_wreq_bits_data_0_ctr; // @[ITTAGE.scala 225:11]
  wire [38:0] table_banks_0_io_wreq_bits_data_0_target; // @[ITTAGE.scala 225:11]
  wire  table_banks_1_clock; // @[ITTAGE.scala 225:11]
  wire  table_banks_1_reset; // @[ITTAGE.scala 225:11]
  wire  table_banks_1_io_rreq_valid; // @[ITTAGE.scala 225:11]
  wire [7:0] table_banks_1_io_rreq_bits_setIdx; // @[ITTAGE.scala 225:11]
  wire [8:0] table_banks_1_io_rresp_data_0_tag; // @[ITTAGE.scala 225:11]
  wire [1:0] table_banks_1_io_rresp_data_0_ctr; // @[ITTAGE.scala 225:11]
  wire [38:0] table_banks_1_io_rresp_data_0_target; // @[ITTAGE.scala 225:11]
  wire  table_banks_1_io_wreq_valid; // @[ITTAGE.scala 225:11]
  wire [7:0] table_banks_1_io_wreq_bits_setIdx; // @[ITTAGE.scala 225:11]
  wire [8:0] table_banks_1_io_wreq_bits_data_0_tag; // @[ITTAGE.scala 225:11]
  wire [1:0] table_banks_1_io_wreq_bits_data_0_ctr; // @[ITTAGE.scala 225:11]
  wire [38:0] table_banks_1_io_wreq_bits_data_0_target; // @[ITTAGE.scala 225:11]
  wire  wrbypass_clock; // @[ITTAGE.scala 276:24]
  wire  wrbypass_reset; // @[ITTAGE.scala 276:24]
  wire  wrbypass_io_wen; // @[ITTAGE.scala 276:24]
  wire [8:0] wrbypass_io_write_idx; // @[ITTAGE.scala 276:24]
  wire [8:0] wrbypass_io_write_tag; // @[ITTAGE.scala 276:24]
  wire [1:0] wrbypass_io_write_data_0; // @[ITTAGE.scala 276:24]
  wire  wrbypass_io_hit; // @[ITTAGE.scala 276:24]
  wire [1:0] wrbypass_io_hit_data_0_bits; // @[ITTAGE.scala 276:24]
  reg [511:0] validArray; // @[ITTAGE.scala 205:27]
  wire [37:0] s0_unhashed_idx = io_req_bits_pc[38:1]; // @[ITTAGE.scala 212:43]
  wire [37:0] _GEN_1031 = {{29'd0}, io_req_bits_folded_hist_hist_7_folded_hist}; // @[ITTAGE.scala 186:31]
  wire [37:0] _idx_T = s0_unhashed_idx ^ _GEN_1031; // @[ITTAGE.scala 186:31]
  wire [8:0] s0_idx = _idx_T[8:0]; // @[ITTAGE.scala 186:40]
  wire [28:0] _GEN_1032 = {{20'd0}, io_req_bits_folded_hist_hist_7_folded_hist}; // @[ITTAGE.scala 187:52]
  wire [28:0] _tag_T_1 = s0_unhashed_idx[37:9] ^ _GEN_1032; // @[ITTAGE.scala 187:52]
  wire [8:0] _tag_T_2 = {io_req_bits_folded_hist_hist_0_folded_hist, 1'h0}; // @[ITTAGE.scala 187:75]
  wire [28:0] _GEN_1033 = {{20'd0}, _tag_T_2}; // @[ITTAGE.scala 187:61]
  wire [28:0] _tag_T_3 = _tag_T_1 ^ _GEN_1033; // @[ITTAGE.scala 187:61]
  wire [8:0] s0_tag = _tag_T_3[8:0]; // @[ITTAGE.scala 187:82]
  wire  _T = io_req_ready & io_req_valid; // @[Decoupled.scala 50:35]
  reg [8:0] s1_idx; // @[Reg.scala 16:16]
  reg [8:0] s1_tag; // @[Reg.scala 16:16]
  wire  s0_bank_req_1h_0 = ~s0_idx[0]; // @[ITTAGE.scala 165:86]
  reg  s1_bank_req_1h_0; // @[Reg.scala 16:16]
  reg  s1_bank_req_1h_1; // @[Reg.scala 16:16]
  wire [38:0] _resp_selected_T = s1_bank_req_1h_0 ? table_banks_0_io_rresp_data_0_target : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _resp_selected_T_1 = s1_bank_req_1h_1 ? table_banks_1_io_rresp_data_0_target : 39'h0; // @[Mux.scala 27:73]
  wire [1:0] _resp_selected_T_3 = s1_bank_req_1h_0 ? table_banks_0_io_rresp_data_0_ctr : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _resp_selected_T_4 = s1_bank_req_1h_1 ? table_banks_1_io_rresp_data_0_ctr : 2'h0; // @[Mux.scala 27:73]
  wire [8:0] _resp_selected_T_6 = s1_bank_req_1h_0 ? table_banks_0_io_rresp_data_0_tag : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _resp_selected_T_7 = s1_bank_req_1h_1 ? table_banks_1_io_rresp_data_0_tag : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] resp_selected_tag = _resp_selected_T_6 | _resp_selected_T_7; // @[Mux.scala 27:73]
  wire [511:0] _s1_req_rhit_T = validArray >> s1_idx; // @[ITTAGE.scala 237:31]
  wire  s1_req_rhit = _s1_req_rhit_T[0] & resp_selected_tag == s1_tag; // @[ITTAGE.scala 237:40]
  reg  s1_bank_has_write_on_this_req_0; // @[Reg.scala 16:16]
  reg  s1_bank_has_write_on_this_req_1; // @[Reg.scala 16:16]
  wire  resp_invalid_by_write = s1_bank_req_1h_0 & s1_bank_has_write_on_this_req_0 | s1_bank_req_1h_1 &
    s1_bank_has_write_on_this_req_1; // @[Mux.scala 27:73]
  wire  _s1_bank_has_write_on_this_req_WIRE_0 = table_banks_0_io_wreq_valid; // @[ITTAGE.scala 245:{56,56}]
  wire  _s1_bank_has_write_on_this_req_WIRE_1 = table_banks_1_io_wreq_valid; // @[ITTAGE.scala 245:{56,56}]
  wire [37:0] _GEN_1034 = {{29'd0}, io_update_folded_hist_hist_7_folded_hist}; // @[ITTAGE.scala 186:31]
  wire [37:0] _idx_T_1 = io_update_pc[38:1] ^ _GEN_1034; // @[ITTAGE.scala 186:31]
  wire [8:0] update_idx = _idx_T_1[8:0]; // @[ITTAGE.scala 186:40]
  wire [28:0] _GEN_1035 = {{20'd0}, io_update_folded_hist_hist_7_folded_hist}; // @[ITTAGE.scala 187:52]
  wire [28:0] _tag_T_5 = io_update_pc[38:10] ^ _GEN_1035; // @[ITTAGE.scala 187:52]
  wire [8:0] _tag_T_6 = {io_update_folded_hist_hist_0_folded_hist, 1'h0}; // @[ITTAGE.scala 187:75]
  wire [28:0] _GEN_1036 = {{20'd0}, _tag_T_6}; // @[ITTAGE.scala 187:61]
  wire [28:0] _tag_T_7 = _tag_T_5 ^ _GEN_1036; // @[ITTAGE.scala 187:61]
  wire  update_req_bank_1h_0 = ~update_idx[0]; // @[ITTAGE.scala 165:86]
  wire [1:0] old_ctr = wrbypass_io_hit ? wrbypass_io_hit_data_0_bits : io_update_oldCtr; // @[ITTAGE.scala 283:20]
  wire  update_wdata_ctr_oldSatTaken = old_ctr == 2'h3; // @[BPU.scala 87:27]
  wire  update_wdata_ctr_oldSatNotTaken = old_ctr == 2'h0; // @[BPU.scala 88:30]
  wire [1:0] _update_wdata_ctr_T_4 = old_ctr + 2'h1; // @[BPU.scala 91:24]
  wire [1:0] _update_wdata_ctr_T_6 = old_ctr - 2'h1; // @[BPU.scala 91:35]
  wire [1:0] _update_wdata_ctr_T_7 = io_update_correct ? _update_wdata_ctr_T_4 : _update_wdata_ctr_T_6; // @[BPU.scala 91:12]
  wire [1:0] _update_wdata_ctr_T_8 = update_wdata_ctr_oldSatNotTaken & ~io_update_correct ? 2'h0 : _update_wdata_ctr_T_7
    ; // @[BPU.scala 90:10]
  wire [1:0] _update_wdata_ctr_T_9 = update_wdata_ctr_oldSatTaken & io_update_correct ? 2'h3 : _update_wdata_ctr_T_8; // @[BPU.scala 89:8]
  wire  _GEN_6 = 9'h0 == update_idx | validArray[0]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_7 = 9'h1 == update_idx | validArray[1]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_8 = 9'h2 == update_idx | validArray[2]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_9 = 9'h3 == update_idx | validArray[3]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_10 = 9'h4 == update_idx | validArray[4]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_11 = 9'h5 == update_idx | validArray[5]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_12 = 9'h6 == update_idx | validArray[6]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_13 = 9'h7 == update_idx | validArray[7]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_14 = 9'h8 == update_idx | validArray[8]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_15 = 9'h9 == update_idx | validArray[9]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_16 = 9'ha == update_idx | validArray[10]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_17 = 9'hb == update_idx | validArray[11]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_18 = 9'hc == update_idx | validArray[12]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_19 = 9'hd == update_idx | validArray[13]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_20 = 9'he == update_idx | validArray[14]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_21 = 9'hf == update_idx | validArray[15]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_22 = 9'h10 == update_idx | validArray[16]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_23 = 9'h11 == update_idx | validArray[17]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_24 = 9'h12 == update_idx | validArray[18]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_25 = 9'h13 == update_idx | validArray[19]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_26 = 9'h14 == update_idx | validArray[20]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_27 = 9'h15 == update_idx | validArray[21]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_28 = 9'h16 == update_idx | validArray[22]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_29 = 9'h17 == update_idx | validArray[23]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_30 = 9'h18 == update_idx | validArray[24]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_31 = 9'h19 == update_idx | validArray[25]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_32 = 9'h1a == update_idx | validArray[26]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_33 = 9'h1b == update_idx | validArray[27]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_34 = 9'h1c == update_idx | validArray[28]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_35 = 9'h1d == update_idx | validArray[29]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_36 = 9'h1e == update_idx | validArray[30]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_37 = 9'h1f == update_idx | validArray[31]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_38 = 9'h20 == update_idx | validArray[32]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_39 = 9'h21 == update_idx | validArray[33]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_40 = 9'h22 == update_idx | validArray[34]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_41 = 9'h23 == update_idx | validArray[35]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_42 = 9'h24 == update_idx | validArray[36]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_43 = 9'h25 == update_idx | validArray[37]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_44 = 9'h26 == update_idx | validArray[38]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_45 = 9'h27 == update_idx | validArray[39]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_46 = 9'h28 == update_idx | validArray[40]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_47 = 9'h29 == update_idx | validArray[41]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_48 = 9'h2a == update_idx | validArray[42]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_49 = 9'h2b == update_idx | validArray[43]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_50 = 9'h2c == update_idx | validArray[44]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_51 = 9'h2d == update_idx | validArray[45]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_52 = 9'h2e == update_idx | validArray[46]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_53 = 9'h2f == update_idx | validArray[47]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_54 = 9'h30 == update_idx | validArray[48]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_55 = 9'h31 == update_idx | validArray[49]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_56 = 9'h32 == update_idx | validArray[50]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_57 = 9'h33 == update_idx | validArray[51]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_58 = 9'h34 == update_idx | validArray[52]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_59 = 9'h35 == update_idx | validArray[53]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_60 = 9'h36 == update_idx | validArray[54]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_61 = 9'h37 == update_idx | validArray[55]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_62 = 9'h38 == update_idx | validArray[56]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_63 = 9'h39 == update_idx | validArray[57]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_64 = 9'h3a == update_idx | validArray[58]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_65 = 9'h3b == update_idx | validArray[59]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_66 = 9'h3c == update_idx | validArray[60]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_67 = 9'h3d == update_idx | validArray[61]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_68 = 9'h3e == update_idx | validArray[62]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_69 = 9'h3f == update_idx | validArray[63]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_70 = 9'h40 == update_idx | validArray[64]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_71 = 9'h41 == update_idx | validArray[65]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_72 = 9'h42 == update_idx | validArray[66]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_73 = 9'h43 == update_idx | validArray[67]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_74 = 9'h44 == update_idx | validArray[68]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_75 = 9'h45 == update_idx | validArray[69]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_76 = 9'h46 == update_idx | validArray[70]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_77 = 9'h47 == update_idx | validArray[71]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_78 = 9'h48 == update_idx | validArray[72]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_79 = 9'h49 == update_idx | validArray[73]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_80 = 9'h4a == update_idx | validArray[74]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_81 = 9'h4b == update_idx | validArray[75]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_82 = 9'h4c == update_idx | validArray[76]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_83 = 9'h4d == update_idx | validArray[77]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_84 = 9'h4e == update_idx | validArray[78]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_85 = 9'h4f == update_idx | validArray[79]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_86 = 9'h50 == update_idx | validArray[80]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_87 = 9'h51 == update_idx | validArray[81]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_88 = 9'h52 == update_idx | validArray[82]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_89 = 9'h53 == update_idx | validArray[83]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_90 = 9'h54 == update_idx | validArray[84]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_91 = 9'h55 == update_idx | validArray[85]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_92 = 9'h56 == update_idx | validArray[86]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_93 = 9'h57 == update_idx | validArray[87]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_94 = 9'h58 == update_idx | validArray[88]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_95 = 9'h59 == update_idx | validArray[89]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_96 = 9'h5a == update_idx | validArray[90]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_97 = 9'h5b == update_idx | validArray[91]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_98 = 9'h5c == update_idx | validArray[92]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_99 = 9'h5d == update_idx | validArray[93]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_100 = 9'h5e == update_idx | validArray[94]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_101 = 9'h5f == update_idx | validArray[95]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_102 = 9'h60 == update_idx | validArray[96]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_103 = 9'h61 == update_idx | validArray[97]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_104 = 9'h62 == update_idx | validArray[98]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_105 = 9'h63 == update_idx | validArray[99]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_106 = 9'h64 == update_idx | validArray[100]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_107 = 9'h65 == update_idx | validArray[101]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_108 = 9'h66 == update_idx | validArray[102]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_109 = 9'h67 == update_idx | validArray[103]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_110 = 9'h68 == update_idx | validArray[104]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_111 = 9'h69 == update_idx | validArray[105]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_112 = 9'h6a == update_idx | validArray[106]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_113 = 9'h6b == update_idx | validArray[107]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_114 = 9'h6c == update_idx | validArray[108]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_115 = 9'h6d == update_idx | validArray[109]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_116 = 9'h6e == update_idx | validArray[110]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_117 = 9'h6f == update_idx | validArray[111]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_118 = 9'h70 == update_idx | validArray[112]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_119 = 9'h71 == update_idx | validArray[113]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_120 = 9'h72 == update_idx | validArray[114]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_121 = 9'h73 == update_idx | validArray[115]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_122 = 9'h74 == update_idx | validArray[116]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_123 = 9'h75 == update_idx | validArray[117]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_124 = 9'h76 == update_idx | validArray[118]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_125 = 9'h77 == update_idx | validArray[119]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_126 = 9'h78 == update_idx | validArray[120]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_127 = 9'h79 == update_idx | validArray[121]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_128 = 9'h7a == update_idx | validArray[122]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_129 = 9'h7b == update_idx | validArray[123]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_130 = 9'h7c == update_idx | validArray[124]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_131 = 9'h7d == update_idx | validArray[125]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_132 = 9'h7e == update_idx | validArray[126]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_133 = 9'h7f == update_idx | validArray[127]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_134 = 9'h80 == update_idx | validArray[128]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_135 = 9'h81 == update_idx | validArray[129]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_136 = 9'h82 == update_idx | validArray[130]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_137 = 9'h83 == update_idx | validArray[131]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_138 = 9'h84 == update_idx | validArray[132]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_139 = 9'h85 == update_idx | validArray[133]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_140 = 9'h86 == update_idx | validArray[134]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_141 = 9'h87 == update_idx | validArray[135]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_142 = 9'h88 == update_idx | validArray[136]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_143 = 9'h89 == update_idx | validArray[137]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_144 = 9'h8a == update_idx | validArray[138]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_145 = 9'h8b == update_idx | validArray[139]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_146 = 9'h8c == update_idx | validArray[140]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_147 = 9'h8d == update_idx | validArray[141]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_148 = 9'h8e == update_idx | validArray[142]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_149 = 9'h8f == update_idx | validArray[143]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_150 = 9'h90 == update_idx | validArray[144]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_151 = 9'h91 == update_idx | validArray[145]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_152 = 9'h92 == update_idx | validArray[146]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_153 = 9'h93 == update_idx | validArray[147]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_154 = 9'h94 == update_idx | validArray[148]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_155 = 9'h95 == update_idx | validArray[149]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_156 = 9'h96 == update_idx | validArray[150]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_157 = 9'h97 == update_idx | validArray[151]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_158 = 9'h98 == update_idx | validArray[152]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_159 = 9'h99 == update_idx | validArray[153]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_160 = 9'h9a == update_idx | validArray[154]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_161 = 9'h9b == update_idx | validArray[155]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_162 = 9'h9c == update_idx | validArray[156]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_163 = 9'h9d == update_idx | validArray[157]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_164 = 9'h9e == update_idx | validArray[158]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_165 = 9'h9f == update_idx | validArray[159]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_166 = 9'ha0 == update_idx | validArray[160]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_167 = 9'ha1 == update_idx | validArray[161]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_168 = 9'ha2 == update_idx | validArray[162]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_169 = 9'ha3 == update_idx | validArray[163]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_170 = 9'ha4 == update_idx | validArray[164]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_171 = 9'ha5 == update_idx | validArray[165]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_172 = 9'ha6 == update_idx | validArray[166]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_173 = 9'ha7 == update_idx | validArray[167]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_174 = 9'ha8 == update_idx | validArray[168]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_175 = 9'ha9 == update_idx | validArray[169]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_176 = 9'haa == update_idx | validArray[170]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_177 = 9'hab == update_idx | validArray[171]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_178 = 9'hac == update_idx | validArray[172]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_179 = 9'had == update_idx | validArray[173]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_180 = 9'hae == update_idx | validArray[174]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_181 = 9'haf == update_idx | validArray[175]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_182 = 9'hb0 == update_idx | validArray[176]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_183 = 9'hb1 == update_idx | validArray[177]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_184 = 9'hb2 == update_idx | validArray[178]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_185 = 9'hb3 == update_idx | validArray[179]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_186 = 9'hb4 == update_idx | validArray[180]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_187 = 9'hb5 == update_idx | validArray[181]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_188 = 9'hb6 == update_idx | validArray[182]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_189 = 9'hb7 == update_idx | validArray[183]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_190 = 9'hb8 == update_idx | validArray[184]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_191 = 9'hb9 == update_idx | validArray[185]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_192 = 9'hba == update_idx | validArray[186]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_193 = 9'hbb == update_idx | validArray[187]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_194 = 9'hbc == update_idx | validArray[188]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_195 = 9'hbd == update_idx | validArray[189]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_196 = 9'hbe == update_idx | validArray[190]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_197 = 9'hbf == update_idx | validArray[191]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_198 = 9'hc0 == update_idx | validArray[192]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_199 = 9'hc1 == update_idx | validArray[193]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_200 = 9'hc2 == update_idx | validArray[194]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_201 = 9'hc3 == update_idx | validArray[195]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_202 = 9'hc4 == update_idx | validArray[196]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_203 = 9'hc5 == update_idx | validArray[197]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_204 = 9'hc6 == update_idx | validArray[198]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_205 = 9'hc7 == update_idx | validArray[199]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_206 = 9'hc8 == update_idx | validArray[200]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_207 = 9'hc9 == update_idx | validArray[201]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_208 = 9'hca == update_idx | validArray[202]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_209 = 9'hcb == update_idx | validArray[203]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_210 = 9'hcc == update_idx | validArray[204]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_211 = 9'hcd == update_idx | validArray[205]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_212 = 9'hce == update_idx | validArray[206]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_213 = 9'hcf == update_idx | validArray[207]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_214 = 9'hd0 == update_idx | validArray[208]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_215 = 9'hd1 == update_idx | validArray[209]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_216 = 9'hd2 == update_idx | validArray[210]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_217 = 9'hd3 == update_idx | validArray[211]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_218 = 9'hd4 == update_idx | validArray[212]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_219 = 9'hd5 == update_idx | validArray[213]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_220 = 9'hd6 == update_idx | validArray[214]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_221 = 9'hd7 == update_idx | validArray[215]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_222 = 9'hd8 == update_idx | validArray[216]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_223 = 9'hd9 == update_idx | validArray[217]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_224 = 9'hda == update_idx | validArray[218]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_225 = 9'hdb == update_idx | validArray[219]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_226 = 9'hdc == update_idx | validArray[220]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_227 = 9'hdd == update_idx | validArray[221]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_228 = 9'hde == update_idx | validArray[222]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_229 = 9'hdf == update_idx | validArray[223]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_230 = 9'he0 == update_idx | validArray[224]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_231 = 9'he1 == update_idx | validArray[225]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_232 = 9'he2 == update_idx | validArray[226]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_233 = 9'he3 == update_idx | validArray[227]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_234 = 9'he4 == update_idx | validArray[228]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_235 = 9'he5 == update_idx | validArray[229]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_236 = 9'he6 == update_idx | validArray[230]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_237 = 9'he7 == update_idx | validArray[231]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_238 = 9'he8 == update_idx | validArray[232]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_239 = 9'he9 == update_idx | validArray[233]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_240 = 9'hea == update_idx | validArray[234]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_241 = 9'heb == update_idx | validArray[235]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_242 = 9'hec == update_idx | validArray[236]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_243 = 9'hed == update_idx | validArray[237]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_244 = 9'hee == update_idx | validArray[238]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_245 = 9'hef == update_idx | validArray[239]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_246 = 9'hf0 == update_idx | validArray[240]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_247 = 9'hf1 == update_idx | validArray[241]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_248 = 9'hf2 == update_idx | validArray[242]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_249 = 9'hf3 == update_idx | validArray[243]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_250 = 9'hf4 == update_idx | validArray[244]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_251 = 9'hf5 == update_idx | validArray[245]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_252 = 9'hf6 == update_idx | validArray[246]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_253 = 9'hf7 == update_idx | validArray[247]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_254 = 9'hf8 == update_idx | validArray[248]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_255 = 9'hf9 == update_idx | validArray[249]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_256 = 9'hfa == update_idx | validArray[250]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_257 = 9'hfb == update_idx | validArray[251]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_258 = 9'hfc == update_idx | validArray[252]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_259 = 9'hfd == update_idx | validArray[253]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_260 = 9'hfe == update_idx | validArray[254]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_261 = 9'hff == update_idx | validArray[255]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_262 = 9'h100 == update_idx | validArray[256]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_263 = 9'h101 == update_idx | validArray[257]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_264 = 9'h102 == update_idx | validArray[258]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_265 = 9'h103 == update_idx | validArray[259]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_266 = 9'h104 == update_idx | validArray[260]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_267 = 9'h105 == update_idx | validArray[261]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_268 = 9'h106 == update_idx | validArray[262]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_269 = 9'h107 == update_idx | validArray[263]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_270 = 9'h108 == update_idx | validArray[264]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_271 = 9'h109 == update_idx | validArray[265]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_272 = 9'h10a == update_idx | validArray[266]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_273 = 9'h10b == update_idx | validArray[267]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_274 = 9'h10c == update_idx | validArray[268]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_275 = 9'h10d == update_idx | validArray[269]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_276 = 9'h10e == update_idx | validArray[270]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_277 = 9'h10f == update_idx | validArray[271]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_278 = 9'h110 == update_idx | validArray[272]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_279 = 9'h111 == update_idx | validArray[273]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_280 = 9'h112 == update_idx | validArray[274]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_281 = 9'h113 == update_idx | validArray[275]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_282 = 9'h114 == update_idx | validArray[276]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_283 = 9'h115 == update_idx | validArray[277]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_284 = 9'h116 == update_idx | validArray[278]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_285 = 9'h117 == update_idx | validArray[279]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_286 = 9'h118 == update_idx | validArray[280]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_287 = 9'h119 == update_idx | validArray[281]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_288 = 9'h11a == update_idx | validArray[282]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_289 = 9'h11b == update_idx | validArray[283]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_290 = 9'h11c == update_idx | validArray[284]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_291 = 9'h11d == update_idx | validArray[285]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_292 = 9'h11e == update_idx | validArray[286]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_293 = 9'h11f == update_idx | validArray[287]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_294 = 9'h120 == update_idx | validArray[288]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_295 = 9'h121 == update_idx | validArray[289]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_296 = 9'h122 == update_idx | validArray[290]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_297 = 9'h123 == update_idx | validArray[291]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_298 = 9'h124 == update_idx | validArray[292]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_299 = 9'h125 == update_idx | validArray[293]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_300 = 9'h126 == update_idx | validArray[294]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_301 = 9'h127 == update_idx | validArray[295]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_302 = 9'h128 == update_idx | validArray[296]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_303 = 9'h129 == update_idx | validArray[297]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_304 = 9'h12a == update_idx | validArray[298]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_305 = 9'h12b == update_idx | validArray[299]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_306 = 9'h12c == update_idx | validArray[300]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_307 = 9'h12d == update_idx | validArray[301]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_308 = 9'h12e == update_idx | validArray[302]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_309 = 9'h12f == update_idx | validArray[303]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_310 = 9'h130 == update_idx | validArray[304]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_311 = 9'h131 == update_idx | validArray[305]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_312 = 9'h132 == update_idx | validArray[306]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_313 = 9'h133 == update_idx | validArray[307]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_314 = 9'h134 == update_idx | validArray[308]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_315 = 9'h135 == update_idx | validArray[309]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_316 = 9'h136 == update_idx | validArray[310]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_317 = 9'h137 == update_idx | validArray[311]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_318 = 9'h138 == update_idx | validArray[312]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_319 = 9'h139 == update_idx | validArray[313]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_320 = 9'h13a == update_idx | validArray[314]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_321 = 9'h13b == update_idx | validArray[315]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_322 = 9'h13c == update_idx | validArray[316]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_323 = 9'h13d == update_idx | validArray[317]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_324 = 9'h13e == update_idx | validArray[318]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_325 = 9'h13f == update_idx | validArray[319]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_326 = 9'h140 == update_idx | validArray[320]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_327 = 9'h141 == update_idx | validArray[321]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_328 = 9'h142 == update_idx | validArray[322]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_329 = 9'h143 == update_idx | validArray[323]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_330 = 9'h144 == update_idx | validArray[324]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_331 = 9'h145 == update_idx | validArray[325]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_332 = 9'h146 == update_idx | validArray[326]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_333 = 9'h147 == update_idx | validArray[327]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_334 = 9'h148 == update_idx | validArray[328]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_335 = 9'h149 == update_idx | validArray[329]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_336 = 9'h14a == update_idx | validArray[330]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_337 = 9'h14b == update_idx | validArray[331]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_338 = 9'h14c == update_idx | validArray[332]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_339 = 9'h14d == update_idx | validArray[333]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_340 = 9'h14e == update_idx | validArray[334]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_341 = 9'h14f == update_idx | validArray[335]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_342 = 9'h150 == update_idx | validArray[336]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_343 = 9'h151 == update_idx | validArray[337]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_344 = 9'h152 == update_idx | validArray[338]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_345 = 9'h153 == update_idx | validArray[339]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_346 = 9'h154 == update_idx | validArray[340]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_347 = 9'h155 == update_idx | validArray[341]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_348 = 9'h156 == update_idx | validArray[342]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_349 = 9'h157 == update_idx | validArray[343]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_350 = 9'h158 == update_idx | validArray[344]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_351 = 9'h159 == update_idx | validArray[345]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_352 = 9'h15a == update_idx | validArray[346]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_353 = 9'h15b == update_idx | validArray[347]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_354 = 9'h15c == update_idx | validArray[348]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_355 = 9'h15d == update_idx | validArray[349]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_356 = 9'h15e == update_idx | validArray[350]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_357 = 9'h15f == update_idx | validArray[351]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_358 = 9'h160 == update_idx | validArray[352]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_359 = 9'h161 == update_idx | validArray[353]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_360 = 9'h162 == update_idx | validArray[354]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_361 = 9'h163 == update_idx | validArray[355]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_362 = 9'h164 == update_idx | validArray[356]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_363 = 9'h165 == update_idx | validArray[357]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_364 = 9'h166 == update_idx | validArray[358]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_365 = 9'h167 == update_idx | validArray[359]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_366 = 9'h168 == update_idx | validArray[360]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_367 = 9'h169 == update_idx | validArray[361]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_368 = 9'h16a == update_idx | validArray[362]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_369 = 9'h16b == update_idx | validArray[363]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_370 = 9'h16c == update_idx | validArray[364]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_371 = 9'h16d == update_idx | validArray[365]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_372 = 9'h16e == update_idx | validArray[366]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_373 = 9'h16f == update_idx | validArray[367]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_374 = 9'h170 == update_idx | validArray[368]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_375 = 9'h171 == update_idx | validArray[369]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_376 = 9'h172 == update_idx | validArray[370]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_377 = 9'h173 == update_idx | validArray[371]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_378 = 9'h174 == update_idx | validArray[372]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_379 = 9'h175 == update_idx | validArray[373]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_380 = 9'h176 == update_idx | validArray[374]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_381 = 9'h177 == update_idx | validArray[375]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_382 = 9'h178 == update_idx | validArray[376]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_383 = 9'h179 == update_idx | validArray[377]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_384 = 9'h17a == update_idx | validArray[378]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_385 = 9'h17b == update_idx | validArray[379]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_386 = 9'h17c == update_idx | validArray[380]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_387 = 9'h17d == update_idx | validArray[381]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_388 = 9'h17e == update_idx | validArray[382]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_389 = 9'h17f == update_idx | validArray[383]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_390 = 9'h180 == update_idx | validArray[384]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_391 = 9'h181 == update_idx | validArray[385]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_392 = 9'h182 == update_idx | validArray[386]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_393 = 9'h183 == update_idx | validArray[387]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_394 = 9'h184 == update_idx | validArray[388]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_395 = 9'h185 == update_idx | validArray[389]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_396 = 9'h186 == update_idx | validArray[390]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_397 = 9'h187 == update_idx | validArray[391]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_398 = 9'h188 == update_idx | validArray[392]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_399 = 9'h189 == update_idx | validArray[393]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_400 = 9'h18a == update_idx | validArray[394]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_401 = 9'h18b == update_idx | validArray[395]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_402 = 9'h18c == update_idx | validArray[396]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_403 = 9'h18d == update_idx | validArray[397]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_404 = 9'h18e == update_idx | validArray[398]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_405 = 9'h18f == update_idx | validArray[399]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_406 = 9'h190 == update_idx | validArray[400]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_407 = 9'h191 == update_idx | validArray[401]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_408 = 9'h192 == update_idx | validArray[402]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_409 = 9'h193 == update_idx | validArray[403]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_410 = 9'h194 == update_idx | validArray[404]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_411 = 9'h195 == update_idx | validArray[405]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_412 = 9'h196 == update_idx | validArray[406]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_413 = 9'h197 == update_idx | validArray[407]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_414 = 9'h198 == update_idx | validArray[408]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_415 = 9'h199 == update_idx | validArray[409]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_416 = 9'h19a == update_idx | validArray[410]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_417 = 9'h19b == update_idx | validArray[411]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_418 = 9'h19c == update_idx | validArray[412]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_419 = 9'h19d == update_idx | validArray[413]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_420 = 9'h19e == update_idx | validArray[414]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_421 = 9'h19f == update_idx | validArray[415]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_422 = 9'h1a0 == update_idx | validArray[416]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_423 = 9'h1a1 == update_idx | validArray[417]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_424 = 9'h1a2 == update_idx | validArray[418]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_425 = 9'h1a3 == update_idx | validArray[419]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_426 = 9'h1a4 == update_idx | validArray[420]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_427 = 9'h1a5 == update_idx | validArray[421]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_428 = 9'h1a6 == update_idx | validArray[422]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_429 = 9'h1a7 == update_idx | validArray[423]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_430 = 9'h1a8 == update_idx | validArray[424]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_431 = 9'h1a9 == update_idx | validArray[425]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_432 = 9'h1aa == update_idx | validArray[426]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_433 = 9'h1ab == update_idx | validArray[427]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_434 = 9'h1ac == update_idx | validArray[428]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_435 = 9'h1ad == update_idx | validArray[429]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_436 = 9'h1ae == update_idx | validArray[430]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_437 = 9'h1af == update_idx | validArray[431]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_438 = 9'h1b0 == update_idx | validArray[432]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_439 = 9'h1b1 == update_idx | validArray[433]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_440 = 9'h1b2 == update_idx | validArray[434]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_441 = 9'h1b3 == update_idx | validArray[435]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_442 = 9'h1b4 == update_idx | validArray[436]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_443 = 9'h1b5 == update_idx | validArray[437]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_444 = 9'h1b6 == update_idx | validArray[438]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_445 = 9'h1b7 == update_idx | validArray[439]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_446 = 9'h1b8 == update_idx | validArray[440]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_447 = 9'h1b9 == update_idx | validArray[441]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_448 = 9'h1ba == update_idx | validArray[442]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_449 = 9'h1bb == update_idx | validArray[443]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_450 = 9'h1bc == update_idx | validArray[444]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_451 = 9'h1bd == update_idx | validArray[445]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_452 = 9'h1be == update_idx | validArray[446]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_453 = 9'h1bf == update_idx | validArray[447]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_454 = 9'h1c0 == update_idx | validArray[448]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_455 = 9'h1c1 == update_idx | validArray[449]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_456 = 9'h1c2 == update_idx | validArray[450]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_457 = 9'h1c3 == update_idx | validArray[451]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_458 = 9'h1c4 == update_idx | validArray[452]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_459 = 9'h1c5 == update_idx | validArray[453]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_460 = 9'h1c6 == update_idx | validArray[454]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_461 = 9'h1c7 == update_idx | validArray[455]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_462 = 9'h1c8 == update_idx | validArray[456]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_463 = 9'h1c9 == update_idx | validArray[457]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_464 = 9'h1ca == update_idx | validArray[458]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_465 = 9'h1cb == update_idx | validArray[459]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_466 = 9'h1cc == update_idx | validArray[460]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_467 = 9'h1cd == update_idx | validArray[461]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_468 = 9'h1ce == update_idx | validArray[462]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_469 = 9'h1cf == update_idx | validArray[463]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_470 = 9'h1d0 == update_idx | validArray[464]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_471 = 9'h1d1 == update_idx | validArray[465]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_472 = 9'h1d2 == update_idx | validArray[466]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_473 = 9'h1d3 == update_idx | validArray[467]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_474 = 9'h1d4 == update_idx | validArray[468]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_475 = 9'h1d5 == update_idx | validArray[469]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_476 = 9'h1d6 == update_idx | validArray[470]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_477 = 9'h1d7 == update_idx | validArray[471]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_478 = 9'h1d8 == update_idx | validArray[472]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_479 = 9'h1d9 == update_idx | validArray[473]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_480 = 9'h1da == update_idx | validArray[474]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_481 = 9'h1db == update_idx | validArray[475]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_482 = 9'h1dc == update_idx | validArray[476]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_483 = 9'h1dd == update_idx | validArray[477]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_484 = 9'h1de == update_idx | validArray[478]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_485 = 9'h1df == update_idx | validArray[479]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_486 = 9'h1e0 == update_idx | validArray[480]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_487 = 9'h1e1 == update_idx | validArray[481]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_488 = 9'h1e2 == update_idx | validArray[482]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_489 = 9'h1e3 == update_idx | validArray[483]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_490 = 9'h1e4 == update_idx | validArray[484]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_491 = 9'h1e5 == update_idx | validArray[485]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_492 = 9'h1e6 == update_idx | validArray[486]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_493 = 9'h1e7 == update_idx | validArray[487]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_494 = 9'h1e8 == update_idx | validArray[488]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_495 = 9'h1e9 == update_idx | validArray[489]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_496 = 9'h1ea == update_idx | validArray[490]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_497 = 9'h1eb == update_idx | validArray[491]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_498 = 9'h1ec == update_idx | validArray[492]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_499 = 9'h1ed == update_idx | validArray[493]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_500 = 9'h1ee == update_idx | validArray[494]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_501 = 9'h1ef == update_idx | validArray[495]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_502 = 9'h1f0 == update_idx | validArray[496]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_503 = 9'h1f1 == update_idx | validArray[497]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_504 = 9'h1f2 == update_idx | validArray[498]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_505 = 9'h1f3 == update_idx | validArray[499]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_506 = 9'h1f4 == update_idx | validArray[500]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_507 = 9'h1f5 == update_idx | validArray[501]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_508 = 9'h1f6 == update_idx | validArray[502]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_509 = 9'h1f7 == update_idx | validArray[503]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_510 = 9'h1f8 == update_idx | validArray[504]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_511 = 9'h1f9 == update_idx | validArray[505]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_512 = 9'h1fa == update_idx | validArray[506]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_513 = 9'h1fb == update_idx | validArray[507]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_514 = 9'h1fc == update_idx | validArray[508]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_515 = 9'h1fd == update_idx | validArray[509]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_516 = 9'h1fe == update_idx | validArray[510]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  _GEN_517 = 9'h1ff == update_idx | validArray[511]; // @[ITTAGE.scala 289:30 291:{31,31}]
  wire  newValidArray_1 = io_update_valid ? _GEN_7 : validArray[1]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_0 = io_update_valid ? _GEN_6 : validArray[0]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_3 = io_update_valid ? _GEN_9 : validArray[3]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_2 = io_update_valid ? _GEN_8 : validArray[2]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_5 = io_update_valid ? _GEN_11 : validArray[5]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_4 = io_update_valid ? _GEN_10 : validArray[4]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_7 = io_update_valid ? _GEN_13 : validArray[7]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_6 = io_update_valid ? _GEN_12 : validArray[6]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_lo_lo_lo_lo_lo = {newValidArray_7,newValidArray_6,newValidArray_5,newValidArray_4,
    newValidArray_3,newValidArray_2,newValidArray_1,newValidArray_0}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_9 = io_update_valid ? _GEN_15 : validArray[9]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_8 = io_update_valid ? _GEN_14 : validArray[8]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_11 = io_update_valid ? _GEN_17 : validArray[11]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_10 = io_update_valid ? _GEN_16 : validArray[10]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_13 = io_update_valid ? _GEN_19 : validArray[13]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_12 = io_update_valid ? _GEN_18 : validArray[12]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_15 = io_update_valid ? _GEN_21 : validArray[15]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_14 = io_update_valid ? _GEN_20 : validArray[14]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_lo_lo_lo_lo_lo = {newValidArray_15,newValidArray_14,newValidArray_13,newValidArray_12,
    newValidArray_11,newValidArray_10,newValidArray_9,newValidArray_8,validArray_lo_lo_lo_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_17 = io_update_valid ? _GEN_23 : validArray[17]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_16 = io_update_valid ? _GEN_22 : validArray[16]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_19 = io_update_valid ? _GEN_25 : validArray[19]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_18 = io_update_valid ? _GEN_24 : validArray[18]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_21 = io_update_valid ? _GEN_27 : validArray[21]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_20 = io_update_valid ? _GEN_26 : validArray[20]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_23 = io_update_valid ? _GEN_29 : validArray[23]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_22 = io_update_valid ? _GEN_28 : validArray[22]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_lo_lo_lo_hi_lo = {newValidArray_23,newValidArray_22,newValidArray_21,newValidArray_20,
    newValidArray_19,newValidArray_18,newValidArray_17,newValidArray_16}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_25 = io_update_valid ? _GEN_31 : validArray[25]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_24 = io_update_valid ? _GEN_30 : validArray[24]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_27 = io_update_valid ? _GEN_33 : validArray[27]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_26 = io_update_valid ? _GEN_32 : validArray[26]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_29 = io_update_valid ? _GEN_35 : validArray[29]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_28 = io_update_valid ? _GEN_34 : validArray[28]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_31 = io_update_valid ? _GEN_37 : validArray[31]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_30 = io_update_valid ? _GEN_36 : validArray[30]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_lo_lo_lo_lo = {newValidArray_31,newValidArray_30,newValidArray_29,newValidArray_28,
    newValidArray_27,newValidArray_26,newValidArray_25,newValidArray_24,validArray_lo_lo_lo_lo_hi_lo,
    validArray_lo_lo_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_33 = io_update_valid ? _GEN_39 : validArray[33]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_32 = io_update_valid ? _GEN_38 : validArray[32]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_35 = io_update_valid ? _GEN_41 : validArray[35]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_34 = io_update_valid ? _GEN_40 : validArray[34]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_37 = io_update_valid ? _GEN_43 : validArray[37]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_36 = io_update_valid ? _GEN_42 : validArray[36]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_39 = io_update_valid ? _GEN_45 : validArray[39]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_38 = io_update_valid ? _GEN_44 : validArray[38]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_lo_lo_hi_lo_lo = {newValidArray_39,newValidArray_38,newValidArray_37,newValidArray_36,
    newValidArray_35,newValidArray_34,newValidArray_33,newValidArray_32}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_41 = io_update_valid ? _GEN_47 : validArray[41]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_40 = io_update_valid ? _GEN_46 : validArray[40]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_43 = io_update_valid ? _GEN_49 : validArray[43]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_42 = io_update_valid ? _GEN_48 : validArray[42]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_45 = io_update_valid ? _GEN_51 : validArray[45]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_44 = io_update_valid ? _GEN_50 : validArray[44]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_47 = io_update_valid ? _GEN_53 : validArray[47]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_46 = io_update_valid ? _GEN_52 : validArray[46]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_lo_lo_lo_hi_lo = {newValidArray_47,newValidArray_46,newValidArray_45,newValidArray_44,
    newValidArray_43,newValidArray_42,newValidArray_41,newValidArray_40,validArray_lo_lo_lo_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_49 = io_update_valid ? _GEN_55 : validArray[49]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_48 = io_update_valid ? _GEN_54 : validArray[48]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_51 = io_update_valid ? _GEN_57 : validArray[51]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_50 = io_update_valid ? _GEN_56 : validArray[50]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_53 = io_update_valid ? _GEN_59 : validArray[53]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_52 = io_update_valid ? _GEN_58 : validArray[52]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_55 = io_update_valid ? _GEN_61 : validArray[55]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_54 = io_update_valid ? _GEN_60 : validArray[54]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_lo_lo_hi_hi_lo = {newValidArray_55,newValidArray_54,newValidArray_53,newValidArray_52,
    newValidArray_51,newValidArray_50,newValidArray_49,newValidArray_48}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_57 = io_update_valid ? _GEN_63 : validArray[57]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_56 = io_update_valid ? _GEN_62 : validArray[56]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_59 = io_update_valid ? _GEN_65 : validArray[59]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_58 = io_update_valid ? _GEN_64 : validArray[58]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_61 = io_update_valid ? _GEN_67 : validArray[61]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_60 = io_update_valid ? _GEN_66 : validArray[60]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_63 = io_update_valid ? _GEN_69 : validArray[63]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_62 = io_update_valid ? _GEN_68 : validArray[62]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_lo_lo_lo_hi = {newValidArray_63,newValidArray_62,newValidArray_61,newValidArray_60,
    newValidArray_59,newValidArray_58,newValidArray_57,newValidArray_56,validArray_lo_lo_lo_hi_hi_lo,
    validArray_lo_lo_lo_hi_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_65 = io_update_valid ? _GEN_71 : validArray[65]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_64 = io_update_valid ? _GEN_70 : validArray[64]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_67 = io_update_valid ? _GEN_73 : validArray[67]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_66 = io_update_valid ? _GEN_72 : validArray[66]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_69 = io_update_valid ? _GEN_75 : validArray[69]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_68 = io_update_valid ? _GEN_74 : validArray[68]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_71 = io_update_valid ? _GEN_77 : validArray[71]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_70 = io_update_valid ? _GEN_76 : validArray[70]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_lo_hi_lo_lo_lo = {newValidArray_71,newValidArray_70,newValidArray_69,newValidArray_68,
    newValidArray_67,newValidArray_66,newValidArray_65,newValidArray_64}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_73 = io_update_valid ? _GEN_79 : validArray[73]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_72 = io_update_valid ? _GEN_78 : validArray[72]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_75 = io_update_valid ? _GEN_81 : validArray[75]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_74 = io_update_valid ? _GEN_80 : validArray[74]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_77 = io_update_valid ? _GEN_83 : validArray[77]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_76 = io_update_valid ? _GEN_82 : validArray[76]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_79 = io_update_valid ? _GEN_85 : validArray[79]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_78 = io_update_valid ? _GEN_84 : validArray[78]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_lo_lo_hi_lo_lo = {newValidArray_79,newValidArray_78,newValidArray_77,newValidArray_76,
    newValidArray_75,newValidArray_74,newValidArray_73,newValidArray_72,validArray_lo_lo_hi_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_81 = io_update_valid ? _GEN_87 : validArray[81]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_80 = io_update_valid ? _GEN_86 : validArray[80]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_83 = io_update_valid ? _GEN_89 : validArray[83]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_82 = io_update_valid ? _GEN_88 : validArray[82]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_85 = io_update_valid ? _GEN_91 : validArray[85]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_84 = io_update_valid ? _GEN_90 : validArray[84]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_87 = io_update_valid ? _GEN_93 : validArray[87]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_86 = io_update_valid ? _GEN_92 : validArray[86]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_lo_hi_lo_hi_lo = {newValidArray_87,newValidArray_86,newValidArray_85,newValidArray_84,
    newValidArray_83,newValidArray_82,newValidArray_81,newValidArray_80}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_89 = io_update_valid ? _GEN_95 : validArray[89]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_88 = io_update_valid ? _GEN_94 : validArray[88]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_91 = io_update_valid ? _GEN_97 : validArray[91]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_90 = io_update_valid ? _GEN_96 : validArray[90]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_93 = io_update_valid ? _GEN_99 : validArray[93]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_92 = io_update_valid ? _GEN_98 : validArray[92]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_95 = io_update_valid ? _GEN_101 : validArray[95]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_94 = io_update_valid ? _GEN_100 : validArray[94]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_lo_lo_hi_lo = {newValidArray_95,newValidArray_94,newValidArray_93,newValidArray_92,
    newValidArray_91,newValidArray_90,newValidArray_89,newValidArray_88,validArray_lo_lo_hi_lo_hi_lo,
    validArray_lo_lo_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_97 = io_update_valid ? _GEN_103 : validArray[97]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_96 = io_update_valid ? _GEN_102 : validArray[96]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_99 = io_update_valid ? _GEN_105 : validArray[99]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_98 = io_update_valid ? _GEN_104 : validArray[98]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_101 = io_update_valid ? _GEN_107 : validArray[101]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_100 = io_update_valid ? _GEN_106 : validArray[100]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_103 = io_update_valid ? _GEN_109 : validArray[103]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_102 = io_update_valid ? _GEN_108 : validArray[102]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_lo_hi_hi_lo_lo = {newValidArray_103,newValidArray_102,newValidArray_101,newValidArray_100,
    newValidArray_99,newValidArray_98,newValidArray_97,newValidArray_96}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_105 = io_update_valid ? _GEN_111 : validArray[105]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_104 = io_update_valid ? _GEN_110 : validArray[104]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_107 = io_update_valid ? _GEN_113 : validArray[107]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_106 = io_update_valid ? _GEN_112 : validArray[106]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_109 = io_update_valid ? _GEN_115 : validArray[109]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_108 = io_update_valid ? _GEN_114 : validArray[108]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_111 = io_update_valid ? _GEN_117 : validArray[111]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_110 = io_update_valid ? _GEN_116 : validArray[110]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_lo_lo_hi_hi_lo = {newValidArray_111,newValidArray_110,newValidArray_109,newValidArray_108,
    newValidArray_107,newValidArray_106,newValidArray_105,newValidArray_104,validArray_lo_lo_hi_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_113 = io_update_valid ? _GEN_119 : validArray[113]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_112 = io_update_valid ? _GEN_118 : validArray[112]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_115 = io_update_valid ? _GEN_121 : validArray[115]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_114 = io_update_valid ? _GEN_120 : validArray[114]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_117 = io_update_valid ? _GEN_123 : validArray[117]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_116 = io_update_valid ? _GEN_122 : validArray[116]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_119 = io_update_valid ? _GEN_125 : validArray[119]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_118 = io_update_valid ? _GEN_124 : validArray[118]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_lo_hi_hi_hi_lo = {newValidArray_119,newValidArray_118,newValidArray_117,newValidArray_116,
    newValidArray_115,newValidArray_114,newValidArray_113,newValidArray_112}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_121 = io_update_valid ? _GEN_127 : validArray[121]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_120 = io_update_valid ? _GEN_126 : validArray[120]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_123 = io_update_valid ? _GEN_129 : validArray[123]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_122 = io_update_valid ? _GEN_128 : validArray[122]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_125 = io_update_valid ? _GEN_131 : validArray[125]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_124 = io_update_valid ? _GEN_130 : validArray[124]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_127 = io_update_valid ? _GEN_133 : validArray[127]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_126 = io_update_valid ? _GEN_132 : validArray[126]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_lo_lo_hi_hi = {newValidArray_127,newValidArray_126,newValidArray_125,newValidArray_124,
    newValidArray_123,newValidArray_122,newValidArray_121,newValidArray_120,validArray_lo_lo_hi_hi_hi_lo,
    validArray_lo_lo_hi_hi_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_129 = io_update_valid ? _GEN_135 : validArray[129]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_128 = io_update_valid ? _GEN_134 : validArray[128]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_131 = io_update_valid ? _GEN_137 : validArray[131]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_130 = io_update_valid ? _GEN_136 : validArray[130]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_133 = io_update_valid ? _GEN_139 : validArray[133]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_132 = io_update_valid ? _GEN_138 : validArray[132]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_135 = io_update_valid ? _GEN_141 : validArray[135]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_134 = io_update_valid ? _GEN_140 : validArray[134]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_hi_lo_lo_lo_lo = {newValidArray_135,newValidArray_134,newValidArray_133,newValidArray_132,
    newValidArray_131,newValidArray_130,newValidArray_129,newValidArray_128}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_137 = io_update_valid ? _GEN_143 : validArray[137]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_136 = io_update_valid ? _GEN_142 : validArray[136]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_139 = io_update_valid ? _GEN_145 : validArray[139]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_138 = io_update_valid ? _GEN_144 : validArray[138]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_141 = io_update_valid ? _GEN_147 : validArray[141]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_140 = io_update_valid ? _GEN_146 : validArray[140]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_143 = io_update_valid ? _GEN_149 : validArray[143]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_142 = io_update_valid ? _GEN_148 : validArray[142]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_lo_hi_lo_lo_lo = {newValidArray_143,newValidArray_142,newValidArray_141,newValidArray_140,
    newValidArray_139,newValidArray_138,newValidArray_137,newValidArray_136,validArray_lo_hi_lo_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_145 = io_update_valid ? _GEN_151 : validArray[145]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_144 = io_update_valid ? _GEN_150 : validArray[144]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_147 = io_update_valid ? _GEN_153 : validArray[147]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_146 = io_update_valid ? _GEN_152 : validArray[146]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_149 = io_update_valid ? _GEN_155 : validArray[149]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_148 = io_update_valid ? _GEN_154 : validArray[148]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_151 = io_update_valid ? _GEN_157 : validArray[151]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_150 = io_update_valid ? _GEN_156 : validArray[150]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_hi_lo_lo_hi_lo = {newValidArray_151,newValidArray_150,newValidArray_149,newValidArray_148,
    newValidArray_147,newValidArray_146,newValidArray_145,newValidArray_144}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_153 = io_update_valid ? _GEN_159 : validArray[153]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_152 = io_update_valid ? _GEN_158 : validArray[152]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_155 = io_update_valid ? _GEN_161 : validArray[155]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_154 = io_update_valid ? _GEN_160 : validArray[154]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_157 = io_update_valid ? _GEN_163 : validArray[157]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_156 = io_update_valid ? _GEN_162 : validArray[156]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_159 = io_update_valid ? _GEN_165 : validArray[159]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_158 = io_update_valid ? _GEN_164 : validArray[158]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_lo_hi_lo_lo = {newValidArray_159,newValidArray_158,newValidArray_157,newValidArray_156,
    newValidArray_155,newValidArray_154,newValidArray_153,newValidArray_152,validArray_lo_hi_lo_lo_hi_lo,
    validArray_lo_hi_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_161 = io_update_valid ? _GEN_167 : validArray[161]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_160 = io_update_valid ? _GEN_166 : validArray[160]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_163 = io_update_valid ? _GEN_169 : validArray[163]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_162 = io_update_valid ? _GEN_168 : validArray[162]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_165 = io_update_valid ? _GEN_171 : validArray[165]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_164 = io_update_valid ? _GEN_170 : validArray[164]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_167 = io_update_valid ? _GEN_173 : validArray[167]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_166 = io_update_valid ? _GEN_172 : validArray[166]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_hi_lo_hi_lo_lo = {newValidArray_167,newValidArray_166,newValidArray_165,newValidArray_164,
    newValidArray_163,newValidArray_162,newValidArray_161,newValidArray_160}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_169 = io_update_valid ? _GEN_175 : validArray[169]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_168 = io_update_valid ? _GEN_174 : validArray[168]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_171 = io_update_valid ? _GEN_177 : validArray[171]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_170 = io_update_valid ? _GEN_176 : validArray[170]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_173 = io_update_valid ? _GEN_179 : validArray[173]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_172 = io_update_valid ? _GEN_178 : validArray[172]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_175 = io_update_valid ? _GEN_181 : validArray[175]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_174 = io_update_valid ? _GEN_180 : validArray[174]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_lo_hi_lo_hi_lo = {newValidArray_175,newValidArray_174,newValidArray_173,newValidArray_172,
    newValidArray_171,newValidArray_170,newValidArray_169,newValidArray_168,validArray_lo_hi_lo_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_177 = io_update_valid ? _GEN_183 : validArray[177]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_176 = io_update_valid ? _GEN_182 : validArray[176]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_179 = io_update_valid ? _GEN_185 : validArray[179]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_178 = io_update_valid ? _GEN_184 : validArray[178]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_181 = io_update_valid ? _GEN_187 : validArray[181]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_180 = io_update_valid ? _GEN_186 : validArray[180]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_183 = io_update_valid ? _GEN_189 : validArray[183]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_182 = io_update_valid ? _GEN_188 : validArray[182]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_hi_lo_hi_hi_lo = {newValidArray_183,newValidArray_182,newValidArray_181,newValidArray_180,
    newValidArray_179,newValidArray_178,newValidArray_177,newValidArray_176}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_185 = io_update_valid ? _GEN_191 : validArray[185]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_184 = io_update_valid ? _GEN_190 : validArray[184]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_187 = io_update_valid ? _GEN_193 : validArray[187]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_186 = io_update_valid ? _GEN_192 : validArray[186]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_189 = io_update_valid ? _GEN_195 : validArray[189]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_188 = io_update_valid ? _GEN_194 : validArray[188]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_191 = io_update_valid ? _GEN_197 : validArray[191]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_190 = io_update_valid ? _GEN_196 : validArray[190]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_lo_hi_lo_hi = {newValidArray_191,newValidArray_190,newValidArray_189,newValidArray_188,
    newValidArray_187,newValidArray_186,newValidArray_185,newValidArray_184,validArray_lo_hi_lo_hi_hi_lo,
    validArray_lo_hi_lo_hi_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_193 = io_update_valid ? _GEN_199 : validArray[193]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_192 = io_update_valid ? _GEN_198 : validArray[192]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_195 = io_update_valid ? _GEN_201 : validArray[195]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_194 = io_update_valid ? _GEN_200 : validArray[194]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_197 = io_update_valid ? _GEN_203 : validArray[197]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_196 = io_update_valid ? _GEN_202 : validArray[196]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_199 = io_update_valid ? _GEN_205 : validArray[199]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_198 = io_update_valid ? _GEN_204 : validArray[198]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_hi_hi_lo_lo_lo = {newValidArray_199,newValidArray_198,newValidArray_197,newValidArray_196,
    newValidArray_195,newValidArray_194,newValidArray_193,newValidArray_192}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_201 = io_update_valid ? _GEN_207 : validArray[201]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_200 = io_update_valid ? _GEN_206 : validArray[200]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_203 = io_update_valid ? _GEN_209 : validArray[203]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_202 = io_update_valid ? _GEN_208 : validArray[202]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_205 = io_update_valid ? _GEN_211 : validArray[205]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_204 = io_update_valid ? _GEN_210 : validArray[204]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_207 = io_update_valid ? _GEN_213 : validArray[207]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_206 = io_update_valid ? _GEN_212 : validArray[206]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_lo_hi_hi_lo_lo = {newValidArray_207,newValidArray_206,newValidArray_205,newValidArray_204,
    newValidArray_203,newValidArray_202,newValidArray_201,newValidArray_200,validArray_lo_hi_hi_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_209 = io_update_valid ? _GEN_215 : validArray[209]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_208 = io_update_valid ? _GEN_214 : validArray[208]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_211 = io_update_valid ? _GEN_217 : validArray[211]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_210 = io_update_valid ? _GEN_216 : validArray[210]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_213 = io_update_valid ? _GEN_219 : validArray[213]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_212 = io_update_valid ? _GEN_218 : validArray[212]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_215 = io_update_valid ? _GEN_221 : validArray[215]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_214 = io_update_valid ? _GEN_220 : validArray[214]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_hi_hi_lo_hi_lo = {newValidArray_215,newValidArray_214,newValidArray_213,newValidArray_212,
    newValidArray_211,newValidArray_210,newValidArray_209,newValidArray_208}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_217 = io_update_valid ? _GEN_223 : validArray[217]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_216 = io_update_valid ? _GEN_222 : validArray[216]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_219 = io_update_valid ? _GEN_225 : validArray[219]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_218 = io_update_valid ? _GEN_224 : validArray[218]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_221 = io_update_valid ? _GEN_227 : validArray[221]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_220 = io_update_valid ? _GEN_226 : validArray[220]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_223 = io_update_valid ? _GEN_229 : validArray[223]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_222 = io_update_valid ? _GEN_228 : validArray[222]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_lo_hi_hi_lo = {newValidArray_223,newValidArray_222,newValidArray_221,newValidArray_220,
    newValidArray_219,newValidArray_218,newValidArray_217,newValidArray_216,validArray_lo_hi_hi_lo_hi_lo,
    validArray_lo_hi_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_225 = io_update_valid ? _GEN_231 : validArray[225]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_224 = io_update_valid ? _GEN_230 : validArray[224]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_227 = io_update_valid ? _GEN_233 : validArray[227]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_226 = io_update_valid ? _GEN_232 : validArray[226]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_229 = io_update_valid ? _GEN_235 : validArray[229]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_228 = io_update_valid ? _GEN_234 : validArray[228]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_231 = io_update_valid ? _GEN_237 : validArray[231]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_230 = io_update_valid ? _GEN_236 : validArray[230]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_hi_hi_hi_lo_lo = {newValidArray_231,newValidArray_230,newValidArray_229,newValidArray_228,
    newValidArray_227,newValidArray_226,newValidArray_225,newValidArray_224}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_233 = io_update_valid ? _GEN_239 : validArray[233]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_232 = io_update_valid ? _GEN_238 : validArray[232]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_235 = io_update_valid ? _GEN_241 : validArray[235]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_234 = io_update_valid ? _GEN_240 : validArray[234]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_237 = io_update_valid ? _GEN_243 : validArray[237]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_236 = io_update_valid ? _GEN_242 : validArray[236]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_239 = io_update_valid ? _GEN_245 : validArray[239]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_238 = io_update_valid ? _GEN_244 : validArray[238]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_lo_hi_hi_hi_lo = {newValidArray_239,newValidArray_238,newValidArray_237,newValidArray_236,
    newValidArray_235,newValidArray_234,newValidArray_233,newValidArray_232,validArray_lo_hi_hi_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_241 = io_update_valid ? _GEN_247 : validArray[241]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_240 = io_update_valid ? _GEN_246 : validArray[240]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_243 = io_update_valid ? _GEN_249 : validArray[243]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_242 = io_update_valid ? _GEN_248 : validArray[242]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_245 = io_update_valid ? _GEN_251 : validArray[245]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_244 = io_update_valid ? _GEN_250 : validArray[244]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_247 = io_update_valid ? _GEN_253 : validArray[247]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_246 = io_update_valid ? _GEN_252 : validArray[246]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_lo_hi_hi_hi_hi_lo = {newValidArray_247,newValidArray_246,newValidArray_245,newValidArray_244,
    newValidArray_243,newValidArray_242,newValidArray_241,newValidArray_240}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_249 = io_update_valid ? _GEN_255 : validArray[249]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_248 = io_update_valid ? _GEN_254 : validArray[248]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_251 = io_update_valid ? _GEN_257 : validArray[251]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_250 = io_update_valid ? _GEN_256 : validArray[250]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_253 = io_update_valid ? _GEN_259 : validArray[253]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_252 = io_update_valid ? _GEN_258 : validArray[252]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_255 = io_update_valid ? _GEN_261 : validArray[255]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_254 = io_update_valid ? _GEN_260 : validArray[254]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_lo_hi_hi_hi = {newValidArray_255,newValidArray_254,newValidArray_253,newValidArray_252,
    newValidArray_251,newValidArray_250,newValidArray_249,newValidArray_248,validArray_lo_hi_hi_hi_hi_lo,
    validArray_lo_hi_hi_hi_lo}; // @[ITTAGE.scala 292:33]
  wire [255:0] validArray_lo = {validArray_lo_hi_hi_hi,validArray_lo_hi_hi_lo,validArray_lo_hi_lo_hi,
    validArray_lo_hi_lo_lo,validArray_lo_lo_hi_hi,validArray_lo_lo_hi_lo,validArray_lo_lo_lo_hi,validArray_lo_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_257 = io_update_valid ? _GEN_263 : validArray[257]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_256 = io_update_valid ? _GEN_262 : validArray[256]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_259 = io_update_valid ? _GEN_265 : validArray[259]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_258 = io_update_valid ? _GEN_264 : validArray[258]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_261 = io_update_valid ? _GEN_267 : validArray[261]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_260 = io_update_valid ? _GEN_266 : validArray[260]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_263 = io_update_valid ? _GEN_269 : validArray[263]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_262 = io_update_valid ? _GEN_268 : validArray[262]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_lo_lo_lo_lo_lo = {newValidArray_263,newValidArray_262,newValidArray_261,newValidArray_260,
    newValidArray_259,newValidArray_258,newValidArray_257,newValidArray_256}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_265 = io_update_valid ? _GEN_271 : validArray[265]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_264 = io_update_valid ? _GEN_270 : validArray[264]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_267 = io_update_valid ? _GEN_273 : validArray[267]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_266 = io_update_valid ? _GEN_272 : validArray[266]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_269 = io_update_valid ? _GEN_275 : validArray[269]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_268 = io_update_valid ? _GEN_274 : validArray[268]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_271 = io_update_valid ? _GEN_277 : validArray[271]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_270 = io_update_valid ? _GEN_276 : validArray[270]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_hi_lo_lo_lo_lo = {newValidArray_271,newValidArray_270,newValidArray_269,newValidArray_268,
    newValidArray_267,newValidArray_266,newValidArray_265,newValidArray_264,validArray_hi_lo_lo_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_273 = io_update_valid ? _GEN_279 : validArray[273]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_272 = io_update_valid ? _GEN_278 : validArray[272]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_275 = io_update_valid ? _GEN_281 : validArray[275]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_274 = io_update_valid ? _GEN_280 : validArray[274]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_277 = io_update_valid ? _GEN_283 : validArray[277]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_276 = io_update_valid ? _GEN_282 : validArray[276]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_279 = io_update_valid ? _GEN_285 : validArray[279]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_278 = io_update_valid ? _GEN_284 : validArray[278]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_lo_lo_lo_hi_lo = {newValidArray_279,newValidArray_278,newValidArray_277,newValidArray_276,
    newValidArray_275,newValidArray_274,newValidArray_273,newValidArray_272}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_281 = io_update_valid ? _GEN_287 : validArray[281]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_280 = io_update_valid ? _GEN_286 : validArray[280]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_283 = io_update_valid ? _GEN_289 : validArray[283]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_282 = io_update_valid ? _GEN_288 : validArray[282]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_285 = io_update_valid ? _GEN_291 : validArray[285]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_284 = io_update_valid ? _GEN_290 : validArray[284]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_287 = io_update_valid ? _GEN_293 : validArray[287]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_286 = io_update_valid ? _GEN_292 : validArray[286]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_hi_lo_lo_lo = {newValidArray_287,newValidArray_286,newValidArray_285,newValidArray_284,
    newValidArray_283,newValidArray_282,newValidArray_281,newValidArray_280,validArray_hi_lo_lo_lo_hi_lo,
    validArray_hi_lo_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_289 = io_update_valid ? _GEN_295 : validArray[289]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_288 = io_update_valid ? _GEN_294 : validArray[288]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_291 = io_update_valid ? _GEN_297 : validArray[291]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_290 = io_update_valid ? _GEN_296 : validArray[290]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_293 = io_update_valid ? _GEN_299 : validArray[293]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_292 = io_update_valid ? _GEN_298 : validArray[292]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_295 = io_update_valid ? _GEN_301 : validArray[295]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_294 = io_update_valid ? _GEN_300 : validArray[294]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_lo_lo_hi_lo_lo = {newValidArray_295,newValidArray_294,newValidArray_293,newValidArray_292,
    newValidArray_291,newValidArray_290,newValidArray_289,newValidArray_288}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_297 = io_update_valid ? _GEN_303 : validArray[297]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_296 = io_update_valid ? _GEN_302 : validArray[296]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_299 = io_update_valid ? _GEN_305 : validArray[299]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_298 = io_update_valid ? _GEN_304 : validArray[298]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_301 = io_update_valid ? _GEN_307 : validArray[301]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_300 = io_update_valid ? _GEN_306 : validArray[300]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_303 = io_update_valid ? _GEN_309 : validArray[303]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_302 = io_update_valid ? _GEN_308 : validArray[302]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_hi_lo_lo_hi_lo = {newValidArray_303,newValidArray_302,newValidArray_301,newValidArray_300,
    newValidArray_299,newValidArray_298,newValidArray_297,newValidArray_296,validArray_hi_lo_lo_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_305 = io_update_valid ? _GEN_311 : validArray[305]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_304 = io_update_valid ? _GEN_310 : validArray[304]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_307 = io_update_valid ? _GEN_313 : validArray[307]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_306 = io_update_valid ? _GEN_312 : validArray[306]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_309 = io_update_valid ? _GEN_315 : validArray[309]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_308 = io_update_valid ? _GEN_314 : validArray[308]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_311 = io_update_valid ? _GEN_317 : validArray[311]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_310 = io_update_valid ? _GEN_316 : validArray[310]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_lo_lo_hi_hi_lo = {newValidArray_311,newValidArray_310,newValidArray_309,newValidArray_308,
    newValidArray_307,newValidArray_306,newValidArray_305,newValidArray_304}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_313 = io_update_valid ? _GEN_319 : validArray[313]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_312 = io_update_valid ? _GEN_318 : validArray[312]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_315 = io_update_valid ? _GEN_321 : validArray[315]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_314 = io_update_valid ? _GEN_320 : validArray[314]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_317 = io_update_valid ? _GEN_323 : validArray[317]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_316 = io_update_valid ? _GEN_322 : validArray[316]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_319 = io_update_valid ? _GEN_325 : validArray[319]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_318 = io_update_valid ? _GEN_324 : validArray[318]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_hi_lo_lo_hi = {newValidArray_319,newValidArray_318,newValidArray_317,newValidArray_316,
    newValidArray_315,newValidArray_314,newValidArray_313,newValidArray_312,validArray_hi_lo_lo_hi_hi_lo,
    validArray_hi_lo_lo_hi_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_321 = io_update_valid ? _GEN_327 : validArray[321]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_320 = io_update_valid ? _GEN_326 : validArray[320]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_323 = io_update_valid ? _GEN_329 : validArray[323]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_322 = io_update_valid ? _GEN_328 : validArray[322]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_325 = io_update_valid ? _GEN_331 : validArray[325]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_324 = io_update_valid ? _GEN_330 : validArray[324]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_327 = io_update_valid ? _GEN_333 : validArray[327]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_326 = io_update_valid ? _GEN_332 : validArray[326]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_lo_hi_lo_lo_lo = {newValidArray_327,newValidArray_326,newValidArray_325,newValidArray_324,
    newValidArray_323,newValidArray_322,newValidArray_321,newValidArray_320}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_329 = io_update_valid ? _GEN_335 : validArray[329]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_328 = io_update_valid ? _GEN_334 : validArray[328]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_331 = io_update_valid ? _GEN_337 : validArray[331]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_330 = io_update_valid ? _GEN_336 : validArray[330]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_333 = io_update_valid ? _GEN_339 : validArray[333]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_332 = io_update_valid ? _GEN_338 : validArray[332]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_335 = io_update_valid ? _GEN_341 : validArray[335]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_334 = io_update_valid ? _GEN_340 : validArray[334]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_hi_lo_hi_lo_lo = {newValidArray_335,newValidArray_334,newValidArray_333,newValidArray_332,
    newValidArray_331,newValidArray_330,newValidArray_329,newValidArray_328,validArray_hi_lo_hi_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_337 = io_update_valid ? _GEN_343 : validArray[337]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_336 = io_update_valid ? _GEN_342 : validArray[336]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_339 = io_update_valid ? _GEN_345 : validArray[339]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_338 = io_update_valid ? _GEN_344 : validArray[338]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_341 = io_update_valid ? _GEN_347 : validArray[341]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_340 = io_update_valid ? _GEN_346 : validArray[340]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_343 = io_update_valid ? _GEN_349 : validArray[343]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_342 = io_update_valid ? _GEN_348 : validArray[342]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_lo_hi_lo_hi_lo = {newValidArray_343,newValidArray_342,newValidArray_341,newValidArray_340,
    newValidArray_339,newValidArray_338,newValidArray_337,newValidArray_336}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_345 = io_update_valid ? _GEN_351 : validArray[345]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_344 = io_update_valid ? _GEN_350 : validArray[344]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_347 = io_update_valid ? _GEN_353 : validArray[347]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_346 = io_update_valid ? _GEN_352 : validArray[346]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_349 = io_update_valid ? _GEN_355 : validArray[349]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_348 = io_update_valid ? _GEN_354 : validArray[348]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_351 = io_update_valid ? _GEN_357 : validArray[351]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_350 = io_update_valid ? _GEN_356 : validArray[350]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_hi_lo_hi_lo = {newValidArray_351,newValidArray_350,newValidArray_349,newValidArray_348,
    newValidArray_347,newValidArray_346,newValidArray_345,newValidArray_344,validArray_hi_lo_hi_lo_hi_lo,
    validArray_hi_lo_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_353 = io_update_valid ? _GEN_359 : validArray[353]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_352 = io_update_valid ? _GEN_358 : validArray[352]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_355 = io_update_valid ? _GEN_361 : validArray[355]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_354 = io_update_valid ? _GEN_360 : validArray[354]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_357 = io_update_valid ? _GEN_363 : validArray[357]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_356 = io_update_valid ? _GEN_362 : validArray[356]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_359 = io_update_valid ? _GEN_365 : validArray[359]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_358 = io_update_valid ? _GEN_364 : validArray[358]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_lo_hi_hi_lo_lo = {newValidArray_359,newValidArray_358,newValidArray_357,newValidArray_356,
    newValidArray_355,newValidArray_354,newValidArray_353,newValidArray_352}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_361 = io_update_valid ? _GEN_367 : validArray[361]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_360 = io_update_valid ? _GEN_366 : validArray[360]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_363 = io_update_valid ? _GEN_369 : validArray[363]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_362 = io_update_valid ? _GEN_368 : validArray[362]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_365 = io_update_valid ? _GEN_371 : validArray[365]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_364 = io_update_valid ? _GEN_370 : validArray[364]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_367 = io_update_valid ? _GEN_373 : validArray[367]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_366 = io_update_valid ? _GEN_372 : validArray[366]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_hi_lo_hi_hi_lo = {newValidArray_367,newValidArray_366,newValidArray_365,newValidArray_364,
    newValidArray_363,newValidArray_362,newValidArray_361,newValidArray_360,validArray_hi_lo_hi_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_369 = io_update_valid ? _GEN_375 : validArray[369]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_368 = io_update_valid ? _GEN_374 : validArray[368]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_371 = io_update_valid ? _GEN_377 : validArray[371]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_370 = io_update_valid ? _GEN_376 : validArray[370]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_373 = io_update_valid ? _GEN_379 : validArray[373]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_372 = io_update_valid ? _GEN_378 : validArray[372]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_375 = io_update_valid ? _GEN_381 : validArray[375]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_374 = io_update_valid ? _GEN_380 : validArray[374]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_lo_hi_hi_hi_lo = {newValidArray_375,newValidArray_374,newValidArray_373,newValidArray_372,
    newValidArray_371,newValidArray_370,newValidArray_369,newValidArray_368}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_377 = io_update_valid ? _GEN_383 : validArray[377]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_376 = io_update_valid ? _GEN_382 : validArray[376]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_379 = io_update_valid ? _GEN_385 : validArray[379]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_378 = io_update_valid ? _GEN_384 : validArray[378]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_381 = io_update_valid ? _GEN_387 : validArray[381]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_380 = io_update_valid ? _GEN_386 : validArray[380]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_383 = io_update_valid ? _GEN_389 : validArray[383]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_382 = io_update_valid ? _GEN_388 : validArray[382]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_hi_lo_hi_hi = {newValidArray_383,newValidArray_382,newValidArray_381,newValidArray_380,
    newValidArray_379,newValidArray_378,newValidArray_377,newValidArray_376,validArray_hi_lo_hi_hi_hi_lo,
    validArray_hi_lo_hi_hi_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_385 = io_update_valid ? _GEN_391 : validArray[385]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_384 = io_update_valid ? _GEN_390 : validArray[384]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_387 = io_update_valid ? _GEN_393 : validArray[387]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_386 = io_update_valid ? _GEN_392 : validArray[386]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_389 = io_update_valid ? _GEN_395 : validArray[389]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_388 = io_update_valid ? _GEN_394 : validArray[388]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_391 = io_update_valid ? _GEN_397 : validArray[391]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_390 = io_update_valid ? _GEN_396 : validArray[390]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_hi_lo_lo_lo_lo = {newValidArray_391,newValidArray_390,newValidArray_389,newValidArray_388,
    newValidArray_387,newValidArray_386,newValidArray_385,newValidArray_384}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_393 = io_update_valid ? _GEN_399 : validArray[393]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_392 = io_update_valid ? _GEN_398 : validArray[392]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_395 = io_update_valid ? _GEN_401 : validArray[395]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_394 = io_update_valid ? _GEN_400 : validArray[394]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_397 = io_update_valid ? _GEN_403 : validArray[397]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_396 = io_update_valid ? _GEN_402 : validArray[396]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_399 = io_update_valid ? _GEN_405 : validArray[399]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_398 = io_update_valid ? _GEN_404 : validArray[398]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_hi_hi_lo_lo_lo = {newValidArray_399,newValidArray_398,newValidArray_397,newValidArray_396,
    newValidArray_395,newValidArray_394,newValidArray_393,newValidArray_392,validArray_hi_hi_lo_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_401 = io_update_valid ? _GEN_407 : validArray[401]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_400 = io_update_valid ? _GEN_406 : validArray[400]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_403 = io_update_valid ? _GEN_409 : validArray[403]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_402 = io_update_valid ? _GEN_408 : validArray[402]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_405 = io_update_valid ? _GEN_411 : validArray[405]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_404 = io_update_valid ? _GEN_410 : validArray[404]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_407 = io_update_valid ? _GEN_413 : validArray[407]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_406 = io_update_valid ? _GEN_412 : validArray[406]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_hi_lo_lo_hi_lo = {newValidArray_407,newValidArray_406,newValidArray_405,newValidArray_404,
    newValidArray_403,newValidArray_402,newValidArray_401,newValidArray_400}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_409 = io_update_valid ? _GEN_415 : validArray[409]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_408 = io_update_valid ? _GEN_414 : validArray[408]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_411 = io_update_valid ? _GEN_417 : validArray[411]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_410 = io_update_valid ? _GEN_416 : validArray[410]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_413 = io_update_valid ? _GEN_419 : validArray[413]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_412 = io_update_valid ? _GEN_418 : validArray[412]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_415 = io_update_valid ? _GEN_421 : validArray[415]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_414 = io_update_valid ? _GEN_420 : validArray[414]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_hi_hi_lo_lo = {newValidArray_415,newValidArray_414,newValidArray_413,newValidArray_412,
    newValidArray_411,newValidArray_410,newValidArray_409,newValidArray_408,validArray_hi_hi_lo_lo_hi_lo,
    validArray_hi_hi_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_417 = io_update_valid ? _GEN_423 : validArray[417]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_416 = io_update_valid ? _GEN_422 : validArray[416]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_419 = io_update_valid ? _GEN_425 : validArray[419]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_418 = io_update_valid ? _GEN_424 : validArray[418]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_421 = io_update_valid ? _GEN_427 : validArray[421]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_420 = io_update_valid ? _GEN_426 : validArray[420]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_423 = io_update_valid ? _GEN_429 : validArray[423]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_422 = io_update_valid ? _GEN_428 : validArray[422]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_hi_lo_hi_lo_lo = {newValidArray_423,newValidArray_422,newValidArray_421,newValidArray_420,
    newValidArray_419,newValidArray_418,newValidArray_417,newValidArray_416}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_425 = io_update_valid ? _GEN_431 : validArray[425]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_424 = io_update_valid ? _GEN_430 : validArray[424]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_427 = io_update_valid ? _GEN_433 : validArray[427]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_426 = io_update_valid ? _GEN_432 : validArray[426]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_429 = io_update_valid ? _GEN_435 : validArray[429]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_428 = io_update_valid ? _GEN_434 : validArray[428]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_431 = io_update_valid ? _GEN_437 : validArray[431]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_430 = io_update_valid ? _GEN_436 : validArray[430]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_hi_hi_lo_hi_lo = {newValidArray_431,newValidArray_430,newValidArray_429,newValidArray_428,
    newValidArray_427,newValidArray_426,newValidArray_425,newValidArray_424,validArray_hi_hi_lo_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_433 = io_update_valid ? _GEN_439 : validArray[433]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_432 = io_update_valid ? _GEN_438 : validArray[432]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_435 = io_update_valid ? _GEN_441 : validArray[435]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_434 = io_update_valid ? _GEN_440 : validArray[434]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_437 = io_update_valid ? _GEN_443 : validArray[437]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_436 = io_update_valid ? _GEN_442 : validArray[436]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_439 = io_update_valid ? _GEN_445 : validArray[439]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_438 = io_update_valid ? _GEN_444 : validArray[438]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_hi_lo_hi_hi_lo = {newValidArray_439,newValidArray_438,newValidArray_437,newValidArray_436,
    newValidArray_435,newValidArray_434,newValidArray_433,newValidArray_432}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_441 = io_update_valid ? _GEN_447 : validArray[441]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_440 = io_update_valid ? _GEN_446 : validArray[440]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_443 = io_update_valid ? _GEN_449 : validArray[443]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_442 = io_update_valid ? _GEN_448 : validArray[442]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_445 = io_update_valid ? _GEN_451 : validArray[445]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_444 = io_update_valid ? _GEN_450 : validArray[444]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_447 = io_update_valid ? _GEN_453 : validArray[447]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_446 = io_update_valid ? _GEN_452 : validArray[446]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_hi_hi_lo_hi = {newValidArray_447,newValidArray_446,newValidArray_445,newValidArray_444,
    newValidArray_443,newValidArray_442,newValidArray_441,newValidArray_440,validArray_hi_hi_lo_hi_hi_lo,
    validArray_hi_hi_lo_hi_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_449 = io_update_valid ? _GEN_455 : validArray[449]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_448 = io_update_valid ? _GEN_454 : validArray[448]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_451 = io_update_valid ? _GEN_457 : validArray[451]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_450 = io_update_valid ? _GEN_456 : validArray[450]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_453 = io_update_valid ? _GEN_459 : validArray[453]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_452 = io_update_valid ? _GEN_458 : validArray[452]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_455 = io_update_valid ? _GEN_461 : validArray[455]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_454 = io_update_valid ? _GEN_460 : validArray[454]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_hi_hi_lo_lo_lo = {newValidArray_455,newValidArray_454,newValidArray_453,newValidArray_452,
    newValidArray_451,newValidArray_450,newValidArray_449,newValidArray_448}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_457 = io_update_valid ? _GEN_463 : validArray[457]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_456 = io_update_valid ? _GEN_462 : validArray[456]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_459 = io_update_valid ? _GEN_465 : validArray[459]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_458 = io_update_valid ? _GEN_464 : validArray[458]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_461 = io_update_valid ? _GEN_467 : validArray[461]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_460 = io_update_valid ? _GEN_466 : validArray[460]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_463 = io_update_valid ? _GEN_469 : validArray[463]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_462 = io_update_valid ? _GEN_468 : validArray[462]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_hi_hi_hi_lo_lo = {newValidArray_463,newValidArray_462,newValidArray_461,newValidArray_460,
    newValidArray_459,newValidArray_458,newValidArray_457,newValidArray_456,validArray_hi_hi_hi_lo_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_465 = io_update_valid ? _GEN_471 : validArray[465]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_464 = io_update_valid ? _GEN_470 : validArray[464]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_467 = io_update_valid ? _GEN_473 : validArray[467]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_466 = io_update_valid ? _GEN_472 : validArray[466]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_469 = io_update_valid ? _GEN_475 : validArray[469]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_468 = io_update_valid ? _GEN_474 : validArray[468]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_471 = io_update_valid ? _GEN_477 : validArray[471]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_470 = io_update_valid ? _GEN_476 : validArray[470]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_hi_hi_lo_hi_lo = {newValidArray_471,newValidArray_470,newValidArray_469,newValidArray_468,
    newValidArray_467,newValidArray_466,newValidArray_465,newValidArray_464}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_473 = io_update_valid ? _GEN_479 : validArray[473]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_472 = io_update_valid ? _GEN_478 : validArray[472]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_475 = io_update_valid ? _GEN_481 : validArray[475]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_474 = io_update_valid ? _GEN_480 : validArray[474]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_477 = io_update_valid ? _GEN_483 : validArray[477]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_476 = io_update_valid ? _GEN_482 : validArray[476]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_479 = io_update_valid ? _GEN_485 : validArray[479]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_478 = io_update_valid ? _GEN_484 : validArray[478]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_hi_hi_hi_lo = {newValidArray_479,newValidArray_478,newValidArray_477,newValidArray_476,
    newValidArray_475,newValidArray_474,newValidArray_473,newValidArray_472,validArray_hi_hi_hi_lo_hi_lo,
    validArray_hi_hi_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_481 = io_update_valid ? _GEN_487 : validArray[481]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_480 = io_update_valid ? _GEN_486 : validArray[480]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_483 = io_update_valid ? _GEN_489 : validArray[483]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_482 = io_update_valid ? _GEN_488 : validArray[482]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_485 = io_update_valid ? _GEN_491 : validArray[485]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_484 = io_update_valid ? _GEN_490 : validArray[484]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_487 = io_update_valid ? _GEN_493 : validArray[487]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_486 = io_update_valid ? _GEN_492 : validArray[486]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_hi_hi_hi_lo_lo = {newValidArray_487,newValidArray_486,newValidArray_485,newValidArray_484,
    newValidArray_483,newValidArray_482,newValidArray_481,newValidArray_480}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_489 = io_update_valid ? _GEN_495 : validArray[489]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_488 = io_update_valid ? _GEN_494 : validArray[488]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_491 = io_update_valid ? _GEN_497 : validArray[491]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_490 = io_update_valid ? _GEN_496 : validArray[490]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_493 = io_update_valid ? _GEN_499 : validArray[493]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_492 = io_update_valid ? _GEN_498 : validArray[492]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_495 = io_update_valid ? _GEN_501 : validArray[495]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_494 = io_update_valid ? _GEN_500 : validArray[494]; // @[ITTAGE.scala 290:26 289:30]
  wire [15:0] validArray_hi_hi_hi_hi_lo = {newValidArray_495,newValidArray_494,newValidArray_493,newValidArray_492,
    newValidArray_491,newValidArray_490,newValidArray_489,newValidArray_488,validArray_hi_hi_hi_hi_lo_lo}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_497 = io_update_valid ? _GEN_503 : validArray[497]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_496 = io_update_valid ? _GEN_502 : validArray[496]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_499 = io_update_valid ? _GEN_505 : validArray[499]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_498 = io_update_valid ? _GEN_504 : validArray[498]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_501 = io_update_valid ? _GEN_507 : validArray[501]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_500 = io_update_valid ? _GEN_506 : validArray[500]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_503 = io_update_valid ? _GEN_509 : validArray[503]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_502 = io_update_valid ? _GEN_508 : validArray[502]; // @[ITTAGE.scala 290:26 289:30]
  wire [7:0] validArray_hi_hi_hi_hi_hi_lo = {newValidArray_503,newValidArray_502,newValidArray_501,newValidArray_500,
    newValidArray_499,newValidArray_498,newValidArray_497,newValidArray_496}; // @[ITTAGE.scala 292:33]
  wire  newValidArray_505 = io_update_valid ? _GEN_511 : validArray[505]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_504 = io_update_valid ? _GEN_510 : validArray[504]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_507 = io_update_valid ? _GEN_513 : validArray[507]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_506 = io_update_valid ? _GEN_512 : validArray[506]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_509 = io_update_valid ? _GEN_515 : validArray[509]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_508 = io_update_valid ? _GEN_514 : validArray[508]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_511 = io_update_valid ? _GEN_517 : validArray[511]; // @[ITTAGE.scala 290:26 289:30]
  wire  newValidArray_510 = io_update_valid ? _GEN_516 : validArray[510]; // @[ITTAGE.scala 290:26 289:30]
  wire [31:0] validArray_hi_hi_hi_hi = {newValidArray_511,newValidArray_510,newValidArray_509,newValidArray_508,
    newValidArray_507,newValidArray_506,newValidArray_505,newValidArray_504,validArray_hi_hi_hi_hi_hi_lo,
    validArray_hi_hi_hi_hi_lo}; // @[ITTAGE.scala 292:33]
  wire [511:0] _validArray_T = {validArray_hi_hi_hi_hi,validArray_hi_hi_hi_lo,validArray_hi_hi_lo_hi,
    validArray_hi_hi_lo_lo,validArray_hi_lo_hi_hi,validArray_hi_lo_hi_lo,validArray_hi_lo_lo_hi,validArray_hi_lo_lo_lo,
    validArray_lo}; // @[ITTAGE.scala 292:33]
  Folded1WDataModuleTemplate_2 us ( // @[ITTAGE.scala 222:18]
    .clock(us_clock),
    .reset(us_reset),
    .io_raddr_0(us_io_raddr_0),
    .io_rdata_0(us_io_rdata_0),
    .io_wen(us_io_wen),
    .io_waddr(us_io_waddr),
    .io_wdata(us_io_wdata),
    .io_resetEn(us_io_resetEn)
  );
  FoldedSRAMTemplate_40 table_banks_0 ( // @[ITTAGE.scala 225:11]
    .clock(table_banks_0_clock),
    .reset(table_banks_0_reset),
    .io_rreq_valid(table_banks_0_io_rreq_valid),
    .io_rreq_bits_setIdx(table_banks_0_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(table_banks_0_io_rresp_data_0_tag),
    .io_rresp_data_0_ctr(table_banks_0_io_rresp_data_0_ctr),
    .io_rresp_data_0_target(table_banks_0_io_rresp_data_0_target),
    .io_wreq_valid(table_banks_0_io_wreq_valid),
    .io_wreq_bits_setIdx(table_banks_0_io_wreq_bits_setIdx),
    .io_wreq_bits_data_0_tag(table_banks_0_io_wreq_bits_data_0_tag),
    .io_wreq_bits_data_0_ctr(table_banks_0_io_wreq_bits_data_0_ctr),
    .io_wreq_bits_data_0_target(table_banks_0_io_wreq_bits_data_0_target)
  );
  FoldedSRAMTemplate_40 table_banks_1 ( // @[ITTAGE.scala 225:11]
    .clock(table_banks_1_clock),
    .reset(table_banks_1_reset),
    .io_rreq_valid(table_banks_1_io_rreq_valid),
    .io_rreq_bits_setIdx(table_banks_1_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(table_banks_1_io_rresp_data_0_tag),
    .io_rresp_data_0_ctr(table_banks_1_io_rresp_data_0_ctr),
    .io_rresp_data_0_target(table_banks_1_io_rresp_data_0_target),
    .io_wreq_valid(table_banks_1_io_wreq_valid),
    .io_wreq_bits_setIdx(table_banks_1_io_wreq_bits_setIdx),
    .io_wreq_bits_data_0_tag(table_banks_1_io_wreq_bits_data_0_tag),
    .io_wreq_bits_data_0_ctr(table_banks_1_io_wreq_bits_data_0_ctr),
    .io_wreq_bits_data_0_target(table_banks_1_io_wreq_bits_data_0_target)
  );
  WrBypass_75 wrbypass ( // @[ITTAGE.scala 276:24]
    .clock(wrbypass_clock),
    .reset(wrbypass_reset),
    .io_wen(wrbypass_io_wen),
    .io_write_idx(wrbypass_io_write_idx),
    .io_write_tag(wrbypass_io_write_tag),
    .io_write_data_0(wrbypass_io_write_data_0),
    .io_hit(wrbypass_io_hit),
    .io_hit_data_0_bits(wrbypass_io_hit_data_0_bits)
  );
  assign io_req_ready = 1'h1; // @[ITTAGE.scala 268:16]
  assign io_resp_valid = s1_req_rhit & ~resp_invalid_by_write; // @[ITTAGE.scala 240:50]
  assign io_resp_bits_ctr = _resp_selected_T_3 | _resp_selected_T_4; // @[Mux.scala 27:73]
  assign io_resp_bits_u = {{1'd0}, us_io_rdata_0}; // @[ITTAGE.scala 242:18]
  assign io_resp_bits_target = _resp_selected_T | _resp_selected_T_1; // @[Mux.scala 27:73]
  assign us_clock = clock;
  assign us_reset = reset;
  assign us_io_raddr_0 = _idx_T[8:0]; // @[ITTAGE.scala 186:40]
  assign us_io_wen = io_update_uValid; // @[ITTAGE.scala 272:13]
  assign us_io_waddr = _idx_T_1[8:0]; // @[ITTAGE.scala 186:40]
  assign us_io_wdata = io_update_u; // @[ITTAGE.scala 274:15]
  assign us_io_resetEn = io_update_reset_u; // @[ITTAGE.scala 296:23]
  assign table_banks_0_clock = clock;
  assign table_banks_0_reset = reset;
  assign table_banks_0_io_rreq_valid = _T & s0_bank_req_1h_0; // @[ITTAGE.scala 228:50]
  assign table_banks_0_io_rreq_bits_setIdx = s0_idx[8:1]; // @[ITTAGE.scala 166:37]
  assign table_banks_0_io_wreq_valid = io_update_valid & update_req_bank_1h_0; // @[ITTAGE.scala 260:33]
  assign table_banks_0_io_wreq_bits_setIdx = update_idx[8:1]; // @[ITTAGE.scala 166:37]
  assign table_banks_0_io_wreq_bits_data_0_tag = _tag_T_7[8:0]; // @[ITTAGE.scala 187:82]
  assign table_banks_0_io_wreq_bits_data_0_ctr = io_update_alloc ? 2'h2 : _update_wdata_ctr_T_9; // @[ITTAGE.scala 284:28]
  assign table_banks_0_io_wreq_bits_data_0_target = io_update_alloc | update_wdata_ctr_oldSatNotTaken ?
    io_update_target : io_update_old_target; // @[ITTAGE.scala 287:29]
  assign table_banks_1_clock = clock;
  assign table_banks_1_reset = reset;
  assign table_banks_1_io_rreq_valid = _T & s0_idx[0]; // @[ITTAGE.scala 228:50]
  assign table_banks_1_io_rreq_bits_setIdx = s0_idx[8:1]; // @[ITTAGE.scala 166:37]
  assign table_banks_1_io_wreq_valid = io_update_valid & update_idx[0]; // @[ITTAGE.scala 260:33]
  assign table_banks_1_io_wreq_bits_setIdx = update_idx[8:1]; // @[ITTAGE.scala 166:37]
  assign table_banks_1_io_wreq_bits_data_0_tag = _tag_T_7[8:0]; // @[ITTAGE.scala 187:82]
  assign table_banks_1_io_wreq_bits_data_0_ctr = io_update_alloc ? 2'h2 : _update_wdata_ctr_T_9; // @[ITTAGE.scala 284:28]
  assign table_banks_1_io_wreq_bits_data_0_target = io_update_alloc | update_wdata_ctr_oldSatNotTaken ?
    io_update_target : io_update_old_target; // @[ITTAGE.scala 287:29]
  assign wrbypass_clock = clock;
  assign wrbypass_reset = reset;
  assign wrbypass_io_wen = io_update_valid; // @[ITTAGE.scala 278:19]
  assign wrbypass_io_write_idx = _idx_T_1[8:0]; // @[ITTAGE.scala 186:40]
  assign wrbypass_io_write_tag = _tag_T_7[8:0]; // @[ITTAGE.scala 187:82]
  assign wrbypass_io_write_data_0 = io_update_alloc ? 2'h2 : _update_wdata_ctr_T_9; // @[ITTAGE.scala 284:28]
  always @(posedge clock) begin
    if (_T) begin // @[Reg.scala 17:18]
      s1_idx <= s0_idx; // @[Reg.scala 17:22]
    end
    if (_T) begin // @[Reg.scala 17:18]
      s1_tag <= s0_tag; // @[Reg.scala 17:22]
    end
    if (_T) begin // @[Reg.scala 17:18]
      s1_bank_req_1h_0 <= s0_bank_req_1h_0; // @[Reg.scala 17:22]
    end
    if (_T) begin // @[Reg.scala 17:18]
      s1_bank_req_1h_1 <= s0_idx[0]; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      s1_bank_has_write_on_this_req_0 <= _s1_bank_has_write_on_this_req_WIRE_0; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      s1_bank_has_write_on_this_req_1 <= _s1_bank_has_write_on_this_req_WIRE_1; // @[Reg.scala 17:22]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ITTAGE.scala 290:26]
      validArray <= 512'h0; // @[ITTAGE.scala 292:16]
    end else if (io_update_valid) begin // @[ITTAGE.scala 205:27]
      validArray <= _validArray_T;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  validArray = _RAND_0[511:0];
  _RAND_1 = {1{`RANDOM}};
  s1_idx = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  s1_tag = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  s1_bank_req_1h_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s1_bank_req_1h_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s1_bank_has_write_on_this_req_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s1_bank_has_write_on_this_req_1 = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    validArray = 512'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

