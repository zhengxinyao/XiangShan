module NegedgeDataModule__8entry_1(
  input         clock,
  input  [2:0]  io_raddr_0,
  output        io_rdata_0_brMask_0,
  output        io_rdata_0_brMask_1,
  output        io_rdata_0_brMask_2,
  output        io_rdata_0_brMask_3,
  output        io_rdata_0_brMask_4,
  output        io_rdata_0_brMask_5,
  output        io_rdata_0_brMask_6,
  output        io_rdata_0_brMask_7,
  output        io_rdata_0_jmpInfo_valid,
  output        io_rdata_0_jmpInfo_bits_0,
  output        io_rdata_0_jmpInfo_bits_1,
  output        io_rdata_0_jmpInfo_bits_2,
  output [2:0]  io_rdata_0_jmpOffset,
  output [38:0] io_rdata_0_jalTarget,
  output        io_rdata_0_rvcMask_0,
  output        io_rdata_0_rvcMask_1,
  output        io_rdata_0_rvcMask_2,
  output        io_rdata_0_rvcMask_3,
  output        io_rdata_0_rvcMask_4,
  output        io_rdata_0_rvcMask_5,
  output        io_rdata_0_rvcMask_6,
  output        io_rdata_0_rvcMask_7,
  input         io_wen_0,
  input  [2:0]  io_waddr_0,
  input         io_wdata_0_brMask_0,
  input         io_wdata_0_brMask_1,
  input         io_wdata_0_brMask_2,
  input         io_wdata_0_brMask_3,
  input         io_wdata_0_brMask_4,
  input         io_wdata_0_brMask_5,
  input         io_wdata_0_brMask_6,
  input         io_wdata_0_brMask_7,
  input         io_wdata_0_jmpInfo_valid,
  input         io_wdata_0_jmpInfo_bits_0,
  input         io_wdata_0_jmpInfo_bits_1,
  input         io_wdata_0_jmpInfo_bits_2,
  input  [2:0]  io_wdata_0_jmpOffset,
  input  [38:0] io_wdata_0_jalTarget,
  input         io_wdata_0_rvcMask_0,
  input         io_wdata_0_rvcMask_1,
  input         io_wdata_0_rvcMask_2,
  input         io_wdata_0_rvcMask_3,
  input         io_wdata_0_rvcMask_4,
  input         io_wdata_0_rvcMask_5,
  input         io_wdata_0_rvcMask_6,
  input         io_wdata_0_rvcMask_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
`endif // RANDOMIZE_REG_INIT
  reg  data_0_brMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_brMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_brMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_brMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_brMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_brMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_brMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_brMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_jmpInfo_valid; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_jmpInfo_bits_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_jmpInfo_bits_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_jmpInfo_bits_2; // @[DataModuleTemplate.scala 168:17]
  reg [2:0] data_0_jmpOffset; // @[DataModuleTemplate.scala 168:17]
  reg [38:0] data_0_jalTarget; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_rvcMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_rvcMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_rvcMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_rvcMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_rvcMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_rvcMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_rvcMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_rvcMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_brMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_brMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_brMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_brMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_brMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_brMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_brMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_brMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_jmpInfo_valid; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_jmpInfo_bits_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_jmpInfo_bits_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_jmpInfo_bits_2; // @[DataModuleTemplate.scala 168:17]
  reg [2:0] data_1_jmpOffset; // @[DataModuleTemplate.scala 168:17]
  reg [38:0] data_1_jalTarget; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_rvcMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_rvcMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_rvcMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_rvcMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_rvcMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_rvcMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_rvcMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_rvcMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_brMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_brMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_brMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_brMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_brMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_brMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_brMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_brMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_jmpInfo_valid; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_jmpInfo_bits_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_jmpInfo_bits_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_jmpInfo_bits_2; // @[DataModuleTemplate.scala 168:17]
  reg [2:0] data_2_jmpOffset; // @[DataModuleTemplate.scala 168:17]
  reg [38:0] data_2_jalTarget; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_rvcMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_rvcMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_rvcMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_rvcMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_rvcMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_rvcMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_rvcMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_rvcMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_brMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_brMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_brMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_brMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_brMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_brMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_brMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_brMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_jmpInfo_valid; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_jmpInfo_bits_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_jmpInfo_bits_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_jmpInfo_bits_2; // @[DataModuleTemplate.scala 168:17]
  reg [2:0] data_3_jmpOffset; // @[DataModuleTemplate.scala 168:17]
  reg [38:0] data_3_jalTarget; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_rvcMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_rvcMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_rvcMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_rvcMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_rvcMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_rvcMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_rvcMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_rvcMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_brMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_brMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_brMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_brMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_brMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_brMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_brMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_brMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_jmpInfo_valid; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_jmpInfo_bits_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_jmpInfo_bits_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_jmpInfo_bits_2; // @[DataModuleTemplate.scala 168:17]
  reg [2:0] data_4_jmpOffset; // @[DataModuleTemplate.scala 168:17]
  reg [38:0] data_4_jalTarget; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_rvcMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_rvcMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_rvcMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_rvcMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_rvcMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_rvcMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_rvcMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_rvcMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_brMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_brMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_brMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_brMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_brMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_brMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_brMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_brMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_jmpInfo_valid; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_jmpInfo_bits_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_jmpInfo_bits_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_jmpInfo_bits_2; // @[DataModuleTemplate.scala 168:17]
  reg [2:0] data_5_jmpOffset; // @[DataModuleTemplate.scala 168:17]
  reg [38:0] data_5_jalTarget; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_rvcMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_rvcMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_rvcMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_rvcMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_rvcMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_rvcMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_rvcMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_rvcMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_brMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_brMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_brMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_brMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_brMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_brMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_brMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_brMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_jmpInfo_valid; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_jmpInfo_bits_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_jmpInfo_bits_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_jmpInfo_bits_2; // @[DataModuleTemplate.scala 168:17]
  reg [2:0] data_6_jmpOffset; // @[DataModuleTemplate.scala 168:17]
  reg [38:0] data_6_jalTarget; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_rvcMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_rvcMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_rvcMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_rvcMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_rvcMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_rvcMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_rvcMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_rvcMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_brMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_brMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_brMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_brMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_brMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_brMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_brMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_brMask_7; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_jmpInfo_valid; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_jmpInfo_bits_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_jmpInfo_bits_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_jmpInfo_bits_2; // @[DataModuleTemplate.scala 168:17]
  reg [2:0] data_7_jmpOffset; // @[DataModuleTemplate.scala 168:17]
  reg [38:0] data_7_jalTarget; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_rvcMask_0; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_rvcMask_1; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_rvcMask_2; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_rvcMask_3; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_rvcMask_4; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_rvcMask_5; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_rvcMask_6; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_rvcMask_7; // @[DataModuleTemplate.scala 168:17]
  wire  read_by_0 = io_wen_0 & io_waddr_0 == io_raddr_0; // @[DataModuleTemplate.scala 176:54]
  wire [7:0] addr_dec = 8'h1 << io_raddr_0; // @[OneHot.scala 64:12]
  wire  _io_rdata_0_T_22 = addr_dec[0] & data_0_rvcMask_0 | addr_dec[1] & data_1_rvcMask_0 | addr_dec[2] &
    data_2_rvcMask_0 | addr_dec[3] & data_3_rvcMask_0 | addr_dec[4] & data_4_rvcMask_0 | addr_dec[5] & data_5_rvcMask_0
     | addr_dec[6] & data_6_rvcMask_0 | addr_dec[7] & data_7_rvcMask_0; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_37 = addr_dec[0] & data_0_rvcMask_1 | addr_dec[1] & data_1_rvcMask_1 | addr_dec[2] &
    data_2_rvcMask_1 | addr_dec[3] & data_3_rvcMask_1 | addr_dec[4] & data_4_rvcMask_1 | addr_dec[5] & data_5_rvcMask_1
     | addr_dec[6] & data_6_rvcMask_1 | addr_dec[7] & data_7_rvcMask_1; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_52 = addr_dec[0] & data_0_rvcMask_2 | addr_dec[1] & data_1_rvcMask_2 | addr_dec[2] &
    data_2_rvcMask_2 | addr_dec[3] & data_3_rvcMask_2 | addr_dec[4] & data_4_rvcMask_2 | addr_dec[5] & data_5_rvcMask_2
     | addr_dec[6] & data_6_rvcMask_2 | addr_dec[7] & data_7_rvcMask_2; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_67 = addr_dec[0] & data_0_rvcMask_3 | addr_dec[1] & data_1_rvcMask_3 | addr_dec[2] &
    data_2_rvcMask_3 | addr_dec[3] & data_3_rvcMask_3 | addr_dec[4] & data_4_rvcMask_3 | addr_dec[5] & data_5_rvcMask_3
     | addr_dec[6] & data_6_rvcMask_3 | addr_dec[7] & data_7_rvcMask_3; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_82 = addr_dec[0] & data_0_rvcMask_4 | addr_dec[1] & data_1_rvcMask_4 | addr_dec[2] &
    data_2_rvcMask_4 | addr_dec[3] & data_3_rvcMask_4 | addr_dec[4] & data_4_rvcMask_4 | addr_dec[5] & data_5_rvcMask_4
     | addr_dec[6] & data_6_rvcMask_4 | addr_dec[7] & data_7_rvcMask_4; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_97 = addr_dec[0] & data_0_rvcMask_5 | addr_dec[1] & data_1_rvcMask_5 | addr_dec[2] &
    data_2_rvcMask_5 | addr_dec[3] & data_3_rvcMask_5 | addr_dec[4] & data_4_rvcMask_5 | addr_dec[5] & data_5_rvcMask_5
     | addr_dec[6] & data_6_rvcMask_5 | addr_dec[7] & data_7_rvcMask_5; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_112 = addr_dec[0] & data_0_rvcMask_6 | addr_dec[1] & data_1_rvcMask_6 | addr_dec[2] &
    data_2_rvcMask_6 | addr_dec[3] & data_3_rvcMask_6 | addr_dec[4] & data_4_rvcMask_6 | addr_dec[5] & data_5_rvcMask_6
     | addr_dec[6] & data_6_rvcMask_6 | addr_dec[7] & data_7_rvcMask_6; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_127 = addr_dec[0] & data_0_rvcMask_7 | addr_dec[1] & data_1_rvcMask_7 | addr_dec[2] &
    data_2_rvcMask_7 | addr_dec[3] & data_3_rvcMask_7 | addr_dec[4] & data_4_rvcMask_7 | addr_dec[5] & data_5_rvcMask_7
     | addr_dec[6] & data_6_rvcMask_7 | addr_dec[7] & data_7_rvcMask_7; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_128 = addr_dec[0] ? data_0_jalTarget : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_129 = addr_dec[1] ? data_1_jalTarget : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_130 = addr_dec[2] ? data_2_jalTarget : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_131 = addr_dec[3] ? data_3_jalTarget : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_132 = addr_dec[4] ? data_4_jalTarget : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_133 = addr_dec[5] ? data_5_jalTarget : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_134 = addr_dec[6] ? data_6_jalTarget : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_135 = addr_dec[7] ? data_7_jalTarget : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_136 = _io_rdata_0_T_128 | _io_rdata_0_T_129; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_137 = _io_rdata_0_T_136 | _io_rdata_0_T_130; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_138 = _io_rdata_0_T_137 | _io_rdata_0_T_131; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_139 = _io_rdata_0_T_138 | _io_rdata_0_T_132; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_140 = _io_rdata_0_T_139 | _io_rdata_0_T_133; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_141 = _io_rdata_0_T_140 | _io_rdata_0_T_134; // @[Mux.scala 27:73]
  wire [38:0] _io_rdata_0_T_142 = _io_rdata_0_T_141 | _io_rdata_0_T_135; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_143 = addr_dec[0] ? data_0_jmpOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_144 = addr_dec[1] ? data_1_jmpOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_145 = addr_dec[2] ? data_2_jmpOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_146 = addr_dec[3] ? data_3_jmpOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_147 = addr_dec[4] ? data_4_jmpOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_148 = addr_dec[5] ? data_5_jmpOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_149 = addr_dec[6] ? data_6_jmpOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_150 = addr_dec[7] ? data_7_jmpOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_151 = _io_rdata_0_T_143 | _io_rdata_0_T_144; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_152 = _io_rdata_0_T_151 | _io_rdata_0_T_145; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_153 = _io_rdata_0_T_152 | _io_rdata_0_T_146; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_154 = _io_rdata_0_T_153 | _io_rdata_0_T_147; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_155 = _io_rdata_0_T_154 | _io_rdata_0_T_148; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_156 = _io_rdata_0_T_155 | _io_rdata_0_T_149; // @[Mux.scala 27:73]
  wire [2:0] _io_rdata_0_T_157 = _io_rdata_0_T_156 | _io_rdata_0_T_150; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_172 = addr_dec[0] & data_0_jmpInfo_bits_0 | addr_dec[1] & data_1_jmpInfo_bits_0 | addr_dec[2] &
    data_2_jmpInfo_bits_0 | addr_dec[3] & data_3_jmpInfo_bits_0 | addr_dec[4] & data_4_jmpInfo_bits_0 | addr_dec[5] &
    data_5_jmpInfo_bits_0 | addr_dec[6] & data_6_jmpInfo_bits_0 | addr_dec[7] & data_7_jmpInfo_bits_0; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_187 = addr_dec[0] & data_0_jmpInfo_bits_1 | addr_dec[1] & data_1_jmpInfo_bits_1 | addr_dec[2] &
    data_2_jmpInfo_bits_1 | addr_dec[3] & data_3_jmpInfo_bits_1 | addr_dec[4] & data_4_jmpInfo_bits_1 | addr_dec[5] &
    data_5_jmpInfo_bits_1 | addr_dec[6] & data_6_jmpInfo_bits_1 | addr_dec[7] & data_7_jmpInfo_bits_1; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_202 = addr_dec[0] & data_0_jmpInfo_bits_2 | addr_dec[1] & data_1_jmpInfo_bits_2 | addr_dec[2] &
    data_2_jmpInfo_bits_2 | addr_dec[3] & data_3_jmpInfo_bits_2 | addr_dec[4] & data_4_jmpInfo_bits_2 | addr_dec[5] &
    data_5_jmpInfo_bits_2 | addr_dec[6] & data_6_jmpInfo_bits_2 | addr_dec[7] & data_7_jmpInfo_bits_2; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_217 = addr_dec[0] & data_0_jmpInfo_valid | addr_dec[1] & data_1_jmpInfo_valid | addr_dec[2] &
    data_2_jmpInfo_valid | addr_dec[3] & data_3_jmpInfo_valid | addr_dec[4] & data_4_jmpInfo_valid | addr_dec[5] &
    data_5_jmpInfo_valid | addr_dec[6] & data_6_jmpInfo_valid | addr_dec[7] & data_7_jmpInfo_valid; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_232 = addr_dec[0] & data_0_brMask_0 | addr_dec[1] & data_1_brMask_0 | addr_dec[2] &
    data_2_brMask_0 | addr_dec[3] & data_3_brMask_0 | addr_dec[4] & data_4_brMask_0 | addr_dec[5] & data_5_brMask_0 |
    addr_dec[6] & data_6_brMask_0 | addr_dec[7] & data_7_brMask_0; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_247 = addr_dec[0] & data_0_brMask_1 | addr_dec[1] & data_1_brMask_1 | addr_dec[2] &
    data_2_brMask_1 | addr_dec[3] & data_3_brMask_1 | addr_dec[4] & data_4_brMask_1 | addr_dec[5] & data_5_brMask_1 |
    addr_dec[6] & data_6_brMask_1 | addr_dec[7] & data_7_brMask_1; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_262 = addr_dec[0] & data_0_brMask_2 | addr_dec[1] & data_1_brMask_2 | addr_dec[2] &
    data_2_brMask_2 | addr_dec[3] & data_3_brMask_2 | addr_dec[4] & data_4_brMask_2 | addr_dec[5] & data_5_brMask_2 |
    addr_dec[6] & data_6_brMask_2 | addr_dec[7] & data_7_brMask_2; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_277 = addr_dec[0] & data_0_brMask_3 | addr_dec[1] & data_1_brMask_3 | addr_dec[2] &
    data_2_brMask_3 | addr_dec[3] & data_3_brMask_3 | addr_dec[4] & data_4_brMask_3 | addr_dec[5] & data_5_brMask_3 |
    addr_dec[6] & data_6_brMask_3 | addr_dec[7] & data_7_brMask_3; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_292 = addr_dec[0] & data_0_brMask_4 | addr_dec[1] & data_1_brMask_4 | addr_dec[2] &
    data_2_brMask_4 | addr_dec[3] & data_3_brMask_4 | addr_dec[4] & data_4_brMask_4 | addr_dec[5] & data_5_brMask_4 |
    addr_dec[6] & data_6_brMask_4 | addr_dec[7] & data_7_brMask_4; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_307 = addr_dec[0] & data_0_brMask_5 | addr_dec[1] & data_1_brMask_5 | addr_dec[2] &
    data_2_brMask_5 | addr_dec[3] & data_3_brMask_5 | addr_dec[4] & data_4_brMask_5 | addr_dec[5] & data_5_brMask_5 |
    addr_dec[6] & data_6_brMask_5 | addr_dec[7] & data_7_brMask_5; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_322 = addr_dec[0] & data_0_brMask_6 | addr_dec[1] & data_1_brMask_6 | addr_dec[2] &
    data_2_brMask_6 | addr_dec[3] & data_3_brMask_6 | addr_dec[4] & data_4_brMask_6 | addr_dec[5] & data_5_brMask_6 |
    addr_dec[6] & data_6_brMask_6 | addr_dec[7] & data_7_brMask_6; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_337 = addr_dec[0] & data_0_brMask_7 | addr_dec[1] & data_1_brMask_7 | addr_dec[2] &
    data_2_brMask_7 | addr_dec[3] & data_3_brMask_7 | addr_dec[4] & data_4_brMask_7 | addr_dec[5] & data_5_brMask_7 |
    addr_dec[6] & data_6_brMask_7 | addr_dec[7] & data_7_brMask_7; // @[Mux.scala 27:73]
  wire [7:0] waddr_dec_0 = 8'h1 << io_waddr_0; // @[OneHot.scala 57:35]
  wire  write_wen_0 = io_wen_0 & waddr_dec_0[0]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_0_1 = io_wen_0 & waddr_dec_0[1]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_0_2 = io_wen_0 & waddr_dec_0[2]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_0_3 = io_wen_0 & waddr_dec_0[3]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_0_4 = io_wen_0 & waddr_dec_0[4]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_0_5 = io_wen_0 & waddr_dec_0[5]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_0_6 = io_wen_0 & waddr_dec_0[6]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_0_7 = io_wen_0 & waddr_dec_0[7]; // @[DataModuleTemplate.scala 188:57]
  assign io_rdata_0_brMask_0 = |read_by_0 ? io_wdata_0_brMask_0 : _io_rdata_0_T_232; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_brMask_1 = |read_by_0 ? io_wdata_0_brMask_1 : _io_rdata_0_T_247; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_brMask_2 = |read_by_0 ? io_wdata_0_brMask_2 : _io_rdata_0_T_262; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_brMask_3 = |read_by_0 ? io_wdata_0_brMask_3 : _io_rdata_0_T_277; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_brMask_4 = |read_by_0 ? io_wdata_0_brMask_4 : _io_rdata_0_T_292; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_brMask_5 = |read_by_0 ? io_wdata_0_brMask_5 : _io_rdata_0_T_307; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_brMask_6 = |read_by_0 ? io_wdata_0_brMask_6 : _io_rdata_0_T_322; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_brMask_7 = |read_by_0 ? io_wdata_0_brMask_7 : _io_rdata_0_T_337; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_jmpInfo_valid = |read_by_0 ? io_wdata_0_jmpInfo_valid : _io_rdata_0_T_217; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_jmpInfo_bits_0 = |read_by_0 ? io_wdata_0_jmpInfo_bits_0 : _io_rdata_0_T_172; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_jmpInfo_bits_1 = |read_by_0 ? io_wdata_0_jmpInfo_bits_1 : _io_rdata_0_T_187; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_jmpInfo_bits_2 = |read_by_0 ? io_wdata_0_jmpInfo_bits_2 : _io_rdata_0_T_202; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_jmpOffset = |read_by_0 ? io_wdata_0_jmpOffset : _io_rdata_0_T_157; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_jalTarget = |read_by_0 ? io_wdata_0_jalTarget : _io_rdata_0_T_142; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_rvcMask_0 = |read_by_0 ? io_wdata_0_rvcMask_0 : _io_rdata_0_T_22; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_rvcMask_1 = |read_by_0 ? io_wdata_0_rvcMask_1 : _io_rdata_0_T_37; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_rvcMask_2 = |read_by_0 ? io_wdata_0_rvcMask_2 : _io_rdata_0_T_52; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_rvcMask_3 = |read_by_0 ? io_wdata_0_rvcMask_3 : _io_rdata_0_T_67; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_rvcMask_4 = |read_by_0 ? io_wdata_0_rvcMask_4 : _io_rdata_0_T_82; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_rvcMask_5 = |read_by_0 ? io_wdata_0_rvcMask_5 : _io_rdata_0_T_97; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_rvcMask_6 = |read_by_0 ? io_wdata_0_rvcMask_6 : _io_rdata_0_T_112; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_rvcMask_7 = |read_by_0 ? io_wdata_0_rvcMask_7 : _io_rdata_0_T_127; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  always @(negedge clock) begin
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_brMask_0 <= io_wdata_0_brMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_brMask_1 <= io_wdata_0_brMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_brMask_2 <= io_wdata_0_brMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_brMask_3 <= io_wdata_0_brMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_brMask_4 <= io_wdata_0_brMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_brMask_5 <= io_wdata_0_brMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_brMask_6 <= io_wdata_0_brMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_brMask_7 <= io_wdata_0_brMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_jmpInfo_valid <= io_wdata_0_jmpInfo_valid; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_jmpInfo_bits_0 <= io_wdata_0_jmpInfo_bits_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_jmpInfo_bits_1 <= io_wdata_0_jmpInfo_bits_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_jmpInfo_bits_2 <= io_wdata_0_jmpInfo_bits_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_jmpOffset <= io_wdata_0_jmpOffset; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_jalTarget <= io_wdata_0_jalTarget; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_rvcMask_0 <= io_wdata_0_rvcMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_rvcMask_1 <= io_wdata_0_rvcMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_rvcMask_2 <= io_wdata_0_rvcMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_rvcMask_3 <= io_wdata_0_rvcMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_rvcMask_4 <= io_wdata_0_rvcMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_rvcMask_5 <= io_wdata_0_rvcMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_rvcMask_6 <= io_wdata_0_rvcMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0) begin // @[DataModuleTemplate.scala 189:42]
      data_0_rvcMask_7 <= io_wdata_0_rvcMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_brMask_0 <= io_wdata_0_brMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_brMask_1 <= io_wdata_0_brMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_brMask_2 <= io_wdata_0_brMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_brMask_3 <= io_wdata_0_brMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_brMask_4 <= io_wdata_0_brMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_brMask_5 <= io_wdata_0_brMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_brMask_6 <= io_wdata_0_brMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_brMask_7 <= io_wdata_0_brMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_jmpInfo_valid <= io_wdata_0_jmpInfo_valid; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_jmpInfo_bits_0 <= io_wdata_0_jmpInfo_bits_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_jmpInfo_bits_1 <= io_wdata_0_jmpInfo_bits_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_jmpInfo_bits_2 <= io_wdata_0_jmpInfo_bits_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_jmpOffset <= io_wdata_0_jmpOffset; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_jalTarget <= io_wdata_0_jalTarget; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_rvcMask_0 <= io_wdata_0_rvcMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_rvcMask_1 <= io_wdata_0_rvcMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_rvcMask_2 <= io_wdata_0_rvcMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_rvcMask_3 <= io_wdata_0_rvcMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_rvcMask_4 <= io_wdata_0_rvcMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_rvcMask_5 <= io_wdata_0_rvcMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_rvcMask_6 <= io_wdata_0_rvcMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_1) begin // @[DataModuleTemplate.scala 189:42]
      data_1_rvcMask_7 <= io_wdata_0_rvcMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_brMask_0 <= io_wdata_0_brMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_brMask_1 <= io_wdata_0_brMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_brMask_2 <= io_wdata_0_brMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_brMask_3 <= io_wdata_0_brMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_brMask_4 <= io_wdata_0_brMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_brMask_5 <= io_wdata_0_brMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_brMask_6 <= io_wdata_0_brMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_brMask_7 <= io_wdata_0_brMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_jmpInfo_valid <= io_wdata_0_jmpInfo_valid; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_jmpInfo_bits_0 <= io_wdata_0_jmpInfo_bits_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_jmpInfo_bits_1 <= io_wdata_0_jmpInfo_bits_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_jmpInfo_bits_2 <= io_wdata_0_jmpInfo_bits_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_jmpOffset <= io_wdata_0_jmpOffset; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_jalTarget <= io_wdata_0_jalTarget; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_rvcMask_0 <= io_wdata_0_rvcMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_rvcMask_1 <= io_wdata_0_rvcMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_rvcMask_2 <= io_wdata_0_rvcMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_rvcMask_3 <= io_wdata_0_rvcMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_rvcMask_4 <= io_wdata_0_rvcMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_rvcMask_5 <= io_wdata_0_rvcMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_rvcMask_6 <= io_wdata_0_rvcMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_2) begin // @[DataModuleTemplate.scala 189:42]
      data_2_rvcMask_7 <= io_wdata_0_rvcMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_brMask_0 <= io_wdata_0_brMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_brMask_1 <= io_wdata_0_brMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_brMask_2 <= io_wdata_0_brMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_brMask_3 <= io_wdata_0_brMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_brMask_4 <= io_wdata_0_brMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_brMask_5 <= io_wdata_0_brMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_brMask_6 <= io_wdata_0_brMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_brMask_7 <= io_wdata_0_brMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_jmpInfo_valid <= io_wdata_0_jmpInfo_valid; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_jmpInfo_bits_0 <= io_wdata_0_jmpInfo_bits_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_jmpInfo_bits_1 <= io_wdata_0_jmpInfo_bits_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_jmpInfo_bits_2 <= io_wdata_0_jmpInfo_bits_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_jmpOffset <= io_wdata_0_jmpOffset; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_jalTarget <= io_wdata_0_jalTarget; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_rvcMask_0 <= io_wdata_0_rvcMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_rvcMask_1 <= io_wdata_0_rvcMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_rvcMask_2 <= io_wdata_0_rvcMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_rvcMask_3 <= io_wdata_0_rvcMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_rvcMask_4 <= io_wdata_0_rvcMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_rvcMask_5 <= io_wdata_0_rvcMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_rvcMask_6 <= io_wdata_0_rvcMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_3) begin // @[DataModuleTemplate.scala 189:42]
      data_3_rvcMask_7 <= io_wdata_0_rvcMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_brMask_0 <= io_wdata_0_brMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_brMask_1 <= io_wdata_0_brMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_brMask_2 <= io_wdata_0_brMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_brMask_3 <= io_wdata_0_brMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_brMask_4 <= io_wdata_0_brMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_brMask_5 <= io_wdata_0_brMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_brMask_6 <= io_wdata_0_brMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_brMask_7 <= io_wdata_0_brMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_jmpInfo_valid <= io_wdata_0_jmpInfo_valid; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_jmpInfo_bits_0 <= io_wdata_0_jmpInfo_bits_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_jmpInfo_bits_1 <= io_wdata_0_jmpInfo_bits_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_jmpInfo_bits_2 <= io_wdata_0_jmpInfo_bits_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_jmpOffset <= io_wdata_0_jmpOffset; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_jalTarget <= io_wdata_0_jalTarget; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_rvcMask_0 <= io_wdata_0_rvcMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_rvcMask_1 <= io_wdata_0_rvcMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_rvcMask_2 <= io_wdata_0_rvcMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_rvcMask_3 <= io_wdata_0_rvcMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_rvcMask_4 <= io_wdata_0_rvcMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_rvcMask_5 <= io_wdata_0_rvcMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_rvcMask_6 <= io_wdata_0_rvcMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_4) begin // @[DataModuleTemplate.scala 189:42]
      data_4_rvcMask_7 <= io_wdata_0_rvcMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_brMask_0 <= io_wdata_0_brMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_brMask_1 <= io_wdata_0_brMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_brMask_2 <= io_wdata_0_brMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_brMask_3 <= io_wdata_0_brMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_brMask_4 <= io_wdata_0_brMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_brMask_5 <= io_wdata_0_brMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_brMask_6 <= io_wdata_0_brMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_brMask_7 <= io_wdata_0_brMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_jmpInfo_valid <= io_wdata_0_jmpInfo_valid; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_jmpInfo_bits_0 <= io_wdata_0_jmpInfo_bits_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_jmpInfo_bits_1 <= io_wdata_0_jmpInfo_bits_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_jmpInfo_bits_2 <= io_wdata_0_jmpInfo_bits_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_jmpOffset <= io_wdata_0_jmpOffset; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_jalTarget <= io_wdata_0_jalTarget; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_rvcMask_0 <= io_wdata_0_rvcMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_rvcMask_1 <= io_wdata_0_rvcMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_rvcMask_2 <= io_wdata_0_rvcMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_rvcMask_3 <= io_wdata_0_rvcMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_rvcMask_4 <= io_wdata_0_rvcMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_rvcMask_5 <= io_wdata_0_rvcMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_rvcMask_6 <= io_wdata_0_rvcMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_5) begin // @[DataModuleTemplate.scala 189:42]
      data_5_rvcMask_7 <= io_wdata_0_rvcMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_brMask_0 <= io_wdata_0_brMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_brMask_1 <= io_wdata_0_brMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_brMask_2 <= io_wdata_0_brMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_brMask_3 <= io_wdata_0_brMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_brMask_4 <= io_wdata_0_brMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_brMask_5 <= io_wdata_0_brMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_brMask_6 <= io_wdata_0_brMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_brMask_7 <= io_wdata_0_brMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_jmpInfo_valid <= io_wdata_0_jmpInfo_valid; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_jmpInfo_bits_0 <= io_wdata_0_jmpInfo_bits_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_jmpInfo_bits_1 <= io_wdata_0_jmpInfo_bits_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_jmpInfo_bits_2 <= io_wdata_0_jmpInfo_bits_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_jmpOffset <= io_wdata_0_jmpOffset; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_jalTarget <= io_wdata_0_jalTarget; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_rvcMask_0 <= io_wdata_0_rvcMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_rvcMask_1 <= io_wdata_0_rvcMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_rvcMask_2 <= io_wdata_0_rvcMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_rvcMask_3 <= io_wdata_0_rvcMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_rvcMask_4 <= io_wdata_0_rvcMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_rvcMask_5 <= io_wdata_0_rvcMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_rvcMask_6 <= io_wdata_0_rvcMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_6) begin // @[DataModuleTemplate.scala 189:42]
      data_6_rvcMask_7 <= io_wdata_0_rvcMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_brMask_0 <= io_wdata_0_brMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_brMask_1 <= io_wdata_0_brMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_brMask_2 <= io_wdata_0_brMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_brMask_3 <= io_wdata_0_brMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_brMask_4 <= io_wdata_0_brMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_brMask_5 <= io_wdata_0_brMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_brMask_6 <= io_wdata_0_brMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_brMask_7 <= io_wdata_0_brMask_7; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_jmpInfo_valid <= io_wdata_0_jmpInfo_valid; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_jmpInfo_bits_0 <= io_wdata_0_jmpInfo_bits_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_jmpInfo_bits_1 <= io_wdata_0_jmpInfo_bits_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_jmpInfo_bits_2 <= io_wdata_0_jmpInfo_bits_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_jmpOffset <= io_wdata_0_jmpOffset; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_jalTarget <= io_wdata_0_jalTarget; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_rvcMask_0 <= io_wdata_0_rvcMask_0; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_rvcMask_1 <= io_wdata_0_rvcMask_1; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_rvcMask_2 <= io_wdata_0_rvcMask_2; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_rvcMask_3 <= io_wdata_0_rvcMask_3; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_rvcMask_4 <= io_wdata_0_rvcMask_4; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_rvcMask_5 <= io_wdata_0_rvcMask_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_rvcMask_6 <= io_wdata_0_rvcMask_6; // @[DataModuleTemplate.scala 190:15]
    end
    if (|write_wen_0_7) begin // @[DataModuleTemplate.scala 189:42]
      data_7_rvcMask_7 <= io_wdata_0_rvcMask_7; // @[DataModuleTemplate.scala 190:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_brMask_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_brMask_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_brMask_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_brMask_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_brMask_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_brMask_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_brMask_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_brMask_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_jmpInfo_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_jmpInfo_bits_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_jmpInfo_bits_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_jmpInfo_bits_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_jmpOffset = _RAND_12[2:0];
  _RAND_13 = {2{`RANDOM}};
  data_0_jalTarget = _RAND_13[38:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_rvcMask_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_rvcMask_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_rvcMask_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_rvcMask_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_rvcMask_4 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_rvcMask_5 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_rvcMask_6 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_rvcMask_7 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  data_1_brMask_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  data_1_brMask_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  data_1_brMask_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  data_1_brMask_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  data_1_brMask_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  data_1_brMask_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  data_1_brMask_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  data_1_brMask_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  data_1_jmpInfo_valid = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  data_1_jmpInfo_bits_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_jmpInfo_bits_1 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_jmpInfo_bits_2 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_jmpOffset = _RAND_34[2:0];
  _RAND_35 = {2{`RANDOM}};
  data_1_jalTarget = _RAND_35[38:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_rvcMask_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_rvcMask_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_rvcMask_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_rvcMask_3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_rvcMask_4 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_rvcMask_5 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_rvcMask_6 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_rvcMask_7 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  data_2_brMask_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  data_2_brMask_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  data_2_brMask_2 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  data_2_brMask_3 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  data_2_brMask_4 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  data_2_brMask_5 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  data_2_brMask_6 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  data_2_brMask_7 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  data_2_jmpInfo_valid = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  data_2_jmpInfo_bits_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  data_2_jmpInfo_bits_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  data_2_jmpInfo_bits_2 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  data_2_jmpOffset = _RAND_56[2:0];
  _RAND_57 = {2{`RANDOM}};
  data_2_jalTarget = _RAND_57[38:0];
  _RAND_58 = {1{`RANDOM}};
  data_2_rvcMask_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  data_2_rvcMask_1 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  data_2_rvcMask_2 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  data_2_rvcMask_3 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  data_2_rvcMask_4 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  data_2_rvcMask_5 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  data_2_rvcMask_6 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  data_2_rvcMask_7 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  data_3_brMask_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  data_3_brMask_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  data_3_brMask_2 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  data_3_brMask_3 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  data_3_brMask_4 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  data_3_brMask_5 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  data_3_brMask_6 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  data_3_brMask_7 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  data_3_jmpInfo_valid = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  data_3_jmpInfo_bits_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  data_3_jmpInfo_bits_1 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  data_3_jmpInfo_bits_2 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  data_3_jmpOffset = _RAND_78[2:0];
  _RAND_79 = {2{`RANDOM}};
  data_3_jalTarget = _RAND_79[38:0];
  _RAND_80 = {1{`RANDOM}};
  data_3_rvcMask_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  data_3_rvcMask_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  data_3_rvcMask_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  data_3_rvcMask_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  data_3_rvcMask_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  data_3_rvcMask_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  data_3_rvcMask_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  data_3_rvcMask_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  data_4_brMask_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  data_4_brMask_1 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  data_4_brMask_2 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  data_4_brMask_3 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  data_4_brMask_4 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  data_4_brMask_5 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  data_4_brMask_6 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  data_4_brMask_7 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  data_4_jmpInfo_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  data_4_jmpInfo_bits_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  data_4_jmpInfo_bits_1 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  data_4_jmpInfo_bits_2 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  data_4_jmpOffset = _RAND_100[2:0];
  _RAND_101 = {2{`RANDOM}};
  data_4_jalTarget = _RAND_101[38:0];
  _RAND_102 = {1{`RANDOM}};
  data_4_rvcMask_0 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  data_4_rvcMask_1 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  data_4_rvcMask_2 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  data_4_rvcMask_3 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  data_4_rvcMask_4 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  data_4_rvcMask_5 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  data_4_rvcMask_6 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  data_4_rvcMask_7 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  data_5_brMask_0 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  data_5_brMask_1 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  data_5_brMask_2 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  data_5_brMask_3 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  data_5_brMask_4 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  data_5_brMask_5 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  data_5_brMask_6 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  data_5_brMask_7 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  data_5_jmpInfo_valid = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  data_5_jmpInfo_bits_0 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  data_5_jmpInfo_bits_1 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  data_5_jmpInfo_bits_2 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  data_5_jmpOffset = _RAND_122[2:0];
  _RAND_123 = {2{`RANDOM}};
  data_5_jalTarget = _RAND_123[38:0];
  _RAND_124 = {1{`RANDOM}};
  data_5_rvcMask_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  data_5_rvcMask_1 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  data_5_rvcMask_2 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  data_5_rvcMask_3 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  data_5_rvcMask_4 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  data_5_rvcMask_5 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  data_5_rvcMask_6 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  data_5_rvcMask_7 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  data_6_brMask_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  data_6_brMask_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  data_6_brMask_2 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  data_6_brMask_3 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  data_6_brMask_4 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  data_6_brMask_5 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  data_6_brMask_6 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  data_6_brMask_7 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  data_6_jmpInfo_valid = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  data_6_jmpInfo_bits_0 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  data_6_jmpInfo_bits_1 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  data_6_jmpInfo_bits_2 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  data_6_jmpOffset = _RAND_144[2:0];
  _RAND_145 = {2{`RANDOM}};
  data_6_jalTarget = _RAND_145[38:0];
  _RAND_146 = {1{`RANDOM}};
  data_6_rvcMask_0 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  data_6_rvcMask_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  data_6_rvcMask_2 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  data_6_rvcMask_3 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  data_6_rvcMask_4 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  data_6_rvcMask_5 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  data_6_rvcMask_6 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  data_6_rvcMask_7 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  data_7_brMask_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  data_7_brMask_1 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  data_7_brMask_2 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  data_7_brMask_3 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  data_7_brMask_4 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  data_7_brMask_5 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  data_7_brMask_6 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  data_7_brMask_7 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  data_7_jmpInfo_valid = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  data_7_jmpInfo_bits_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  data_7_jmpInfo_bits_1 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  data_7_jmpInfo_bits_2 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  data_7_jmpOffset = _RAND_166[2:0];
  _RAND_167 = {2{`RANDOM}};
  data_7_jalTarget = _RAND_167[38:0];
  _RAND_168 = {1{`RANDOM}};
  data_7_rvcMask_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  data_7_rvcMask_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  data_7_rvcMask_2 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  data_7_rvcMask_3 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  data_7_rvcMask_4 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  data_7_rvcMask_5 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  data_7_rvcMask_6 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  data_7_rvcMask_7 = _RAND_175[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

