module AXI4Deinterleaver(
  input          clock,
  input          reset,
  output         auto_in_awready,
  input          auto_in_awvalid,
  input  [5:0]   auto_in_awid,
  input  [35:0]  auto_in_awaddr,
  input  [7:0]   auto_in_awlen,
  input  [2:0]   auto_in_awsize,
  input  [1:0]   auto_in_awburst,
  input          auto_in_awlock,
  input  [3:0]   auto_in_awcache,
  input  [2:0]   auto_in_awprot,
  input  [3:0]   auto_in_awqos,
  input  [3:0]   auto_in_awecho_tl_state_size,
  input  [5:0]   auto_in_awecho_tl_state_source,
  output         auto_in_wready,
  input          auto_in_wvalid,
  input  [255:0] auto_in_wdata,
  input  [31:0]  auto_in_wstrb,
  input          auto_in_wlast,
  input          auto_in_bready,
  output         auto_in_bvalid,
  output [5:0]   auto_in_bid,
  output [1:0]   auto_in_bresp,
  output [3:0]   auto_in_becho_tl_state_size,
  output [5:0]   auto_in_becho_tl_state_source,
  output         auto_in_arready,
  input          auto_in_arvalid,
  input  [5:0]   auto_in_arid,
  input  [35:0]  auto_in_araddr,
  input  [7:0]   auto_in_arlen,
  input  [2:0]   auto_in_arsize,
  input  [1:0]   auto_in_arburst,
  input          auto_in_arlock,
  input  [3:0]   auto_in_arcache,
  input  [2:0]   auto_in_arprot,
  input  [3:0]   auto_in_arqos,
  input  [3:0]   auto_in_arecho_tl_state_size,
  input  [5:0]   auto_in_arecho_tl_state_source,
  input          auto_in_rready,
  output         auto_in_rvalid,
  output [5:0]   auto_in_rid,
  output [255:0] auto_in_rdata,
  output [1:0]   auto_in_rresp,
  output [3:0]   auto_in_recho_tl_state_size,
  output [5:0]   auto_in_recho_tl_state_source,
  output         auto_in_rlast,
  input          auto_out_awready,
  output         auto_out_awvalid,
  output [5:0]   auto_out_awid,
  output [35:0]  auto_out_awaddr,
  output [7:0]   auto_out_awlen,
  output [2:0]   auto_out_awsize,
  output [1:0]   auto_out_awburst,
  output         auto_out_awlock,
  output [3:0]   auto_out_awcache,
  output [2:0]   auto_out_awprot,
  output [3:0]   auto_out_awqos,
  output [3:0]   auto_out_awecho_tl_state_size,
  output [5:0]   auto_out_awecho_tl_state_source,
  input          auto_out_wready,
  output         auto_out_wvalid,
  output [255:0] auto_out_wdata,
  output [31:0]  auto_out_wstrb,
  output         auto_out_wlast,
  output         auto_out_bready,
  input          auto_out_bvalid,
  input  [5:0]   auto_out_bid,
  input  [1:0]   auto_out_bresp,
  input  [3:0]   auto_out_becho_tl_state_size,
  input  [5:0]   auto_out_becho_tl_state_source,
  input          auto_out_arready,
  output         auto_out_arvalid,
  output [5:0]   auto_out_arid,
  output [35:0]  auto_out_araddr,
  output [7:0]   auto_out_arlen,
  output [2:0]   auto_out_arsize,
  output [1:0]   auto_out_arburst,
  output         auto_out_arlock,
  output [3:0]   auto_out_arcache,
  output [2:0]   auto_out_arprot,
  output [3:0]   auto_out_arqos,
  output [3:0]   auto_out_arecho_tl_state_size,
  output [5:0]   auto_out_arecho_tl_state_source,
  output         auto_out_rready,
  input          auto_out_rvalid,
  input  [5:0]   auto_out_rid,
  input  [255:0] auto_out_rdata,
  input  [1:0]   auto_out_rresp,
  input  [3:0]   auto_out_recho_tl_state_size,
  input  [5:0]   auto_out_recho_tl_state_source,
  input          auto_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  wire  qs_queue_0_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_0_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_0_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_0_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_0_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_0_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_0_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_0_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_0_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_0_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_0_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_0_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_0_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_0_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_0_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_0_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_0_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_0_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_1_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_1_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_1_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_1_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_1_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_1_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_1_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_1_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_1_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_1_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_1_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_1_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_1_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_1_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_1_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_1_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_1_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_1_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_2_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_2_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_2_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_2_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_2_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_2_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_2_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_2_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_2_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_2_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_2_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_2_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_2_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_2_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_2_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_2_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_2_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_2_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_3_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_3_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_3_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_3_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_3_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_3_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_3_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_3_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_3_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_3_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_3_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_3_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_3_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_3_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_3_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_3_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_3_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_3_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_4_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_4_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_4_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_4_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_4_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_4_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_4_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_4_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_4_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_4_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_4_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_4_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_4_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_4_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_4_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_4_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_4_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_4_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_5_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_5_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_5_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_5_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_5_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_5_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_5_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_5_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_5_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_5_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_5_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_5_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_5_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_5_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_5_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_5_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_5_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_5_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_6_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_6_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_6_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_6_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_6_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_6_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_6_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_6_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_6_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_6_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_6_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_6_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_6_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_6_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_6_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_6_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_6_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_6_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_7_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_7_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_7_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_7_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_7_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_7_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_7_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_7_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_7_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_7_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_7_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_7_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_7_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_7_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_7_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_7_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_7_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_7_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_8_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_8_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_8_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_8_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_8_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_8_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_8_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_8_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_8_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_8_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_8_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_8_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_8_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_8_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_8_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_8_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_8_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_8_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_9_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_9_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_9_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_9_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_9_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_9_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_9_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_9_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_9_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_9_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_9_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_9_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_9_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_9_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_9_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_9_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_9_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_9_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_10_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_10_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_10_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_10_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_10_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_10_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_10_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_10_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_10_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_10_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_10_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_10_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_10_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_10_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_10_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_10_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_10_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_10_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_11_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_11_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_11_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_11_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_11_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_11_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_11_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_11_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_11_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_11_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_11_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_11_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_11_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_11_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_11_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_11_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_11_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_11_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_12_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_12_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_12_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_12_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_12_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_12_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_12_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_12_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_12_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_12_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_12_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_12_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_12_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_12_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_12_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_12_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_12_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_12_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_13_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_13_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_13_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_13_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_13_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_13_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_13_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_13_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_13_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_13_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_13_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_13_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_13_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_13_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_13_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_13_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_13_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_13_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_14_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_14_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_14_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_14_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_14_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_14_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_14_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_14_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_14_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_14_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_14_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_14_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_14_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_14_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_14_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_14_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_14_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_14_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_15_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_15_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_15_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_15_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_15_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_15_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_15_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_15_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_15_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_15_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_15_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_15_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_15_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_15_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_15_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_15_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_15_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_15_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_16_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_16_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_16_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_16_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_16_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_16_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_16_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_16_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_16_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_16_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_16_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_16_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_16_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_16_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_16_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_16_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_16_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_16_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_17_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_17_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_17_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_17_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_17_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_17_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_17_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_17_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_17_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_17_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_17_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_17_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_17_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_17_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_17_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_17_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_17_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_17_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_18_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_18_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_18_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_18_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_18_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_18_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_18_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_18_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_18_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_18_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_18_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_18_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_18_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_18_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_18_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_18_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_18_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_18_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_19_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_19_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_19_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_19_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_19_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_19_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_19_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_19_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_19_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_19_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_19_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_19_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_19_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_19_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_19_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_19_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_19_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_19_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_20_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_20_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_20_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_20_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_20_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_20_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_20_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_20_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_20_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_20_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_20_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_20_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_20_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_20_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_20_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_20_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_20_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_20_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_21_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_21_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_21_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_21_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_21_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_21_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_21_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_21_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_21_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_21_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_21_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_21_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_21_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_21_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_21_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_21_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_21_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_21_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_22_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_22_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_22_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_22_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_22_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_22_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_22_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_22_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_22_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_22_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_22_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_22_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_22_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_22_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_22_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_22_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_22_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_22_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_23_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_23_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_23_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_23_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_23_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_23_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_23_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_23_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_23_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_23_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_23_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_23_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_23_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_23_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_23_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_23_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_23_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_23_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_24_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_24_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_24_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_24_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_24_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_24_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_24_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_24_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_24_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_24_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_24_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_24_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_24_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_24_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_24_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_24_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_24_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_24_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_25_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_25_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_25_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_25_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_25_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_25_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_25_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_25_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_25_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_25_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_25_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_25_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_25_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_25_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_25_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_25_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_25_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_25_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_26_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_26_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_26_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_26_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_26_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_26_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_26_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_26_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_26_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_26_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_26_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_26_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_26_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_26_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_26_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_26_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_26_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_26_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_27_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_27_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_27_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_27_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_27_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_27_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_27_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_27_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_27_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_27_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_27_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_27_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_27_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_27_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_27_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_27_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_27_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_27_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_28_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_28_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_28_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_28_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_28_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_28_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_28_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_28_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_28_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_28_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_28_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_28_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_28_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_28_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_28_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_28_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_28_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_28_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_29_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_29_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_29_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_29_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_29_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_29_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_29_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_29_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_29_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_29_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_29_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_29_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_29_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_29_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_29_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_29_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_29_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_29_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_30_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_30_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_30_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_30_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_30_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_30_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_30_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_30_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_30_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_30_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_30_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_30_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_30_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_30_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_30_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_30_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_30_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_30_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_31_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_31_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_31_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_31_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_31_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_31_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_31_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_31_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_31_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_31_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_31_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_31_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_31_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_31_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_31_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_31_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_31_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_31_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_32_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_32_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_32_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_32_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_32_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_32_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_32_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_32_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_32_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_32_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_32_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_32_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_32_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_32_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_32_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_32_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_32_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_32_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_33_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_33_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_33_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_33_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_33_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_33_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_33_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_33_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_33_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_33_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_33_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_33_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_33_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_33_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_33_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_33_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_33_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_33_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_34_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_34_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_34_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_34_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_34_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_34_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_34_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_34_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_34_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_34_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_34_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_34_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_34_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_34_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_34_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_34_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_34_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_34_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_35_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_35_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_35_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_35_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_35_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_35_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_35_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_35_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_35_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_35_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_35_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_35_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_35_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_35_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_35_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_35_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_35_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_35_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_36_clock; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_36_reset; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_36_io_enq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_36_io_enq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_36_io_enq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_36_io_enq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_36_io_enq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_36_io_enq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_36_io_enq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_36_io_enq_bits_last; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_36_io_deq_ready; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_36_io_deq_valid; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_36_io_deq_bits_id; // @[Deinterleaver.scala 66:27]
  wire [255:0] qs_queue_36_io_deq_bits_data; // @[Deinterleaver.scala 66:27]
  wire [1:0] qs_queue_36_io_deq_bits_resp; // @[Deinterleaver.scala 66:27]
  wire [3:0] qs_queue_36_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 66:27]
  wire [5:0] qs_queue_36_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 66:27]
  wire  qs_queue_36_io_deq_bits_last; // @[Deinterleaver.scala 66:27]
  reg  locked; // @[Deinterleaver.scala 82:29]
  reg [5:0] deq_id; // @[Deinterleaver.scala 83:25]
  wire [63:0] _deq_OH_T = 64'h1 << deq_id; // @[OneHot.scala 64:12]
  wire [36:0] deq_OH = _deq_OH_T[36:0]; // @[OneHot.scala 64:27]
  wire [63:0] _enq_OH_T = 64'h1 << auto_out_rid; // @[OneHot.scala 64:12]
  wire [36:0] enq_OH = _enq_OH_T[36:0]; // @[OneHot.scala 64:27]
  reg [1:0] pending_count; // @[Deinterleaver.scala 92:32]
  wire  enq_readys_36 = qs_queue_36_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_35 = qs_queue_35_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_34 = qs_queue_34_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_33 = qs_queue_33_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_32 = qs_queue_32_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_31 = qs_queue_31_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_30 = qs_queue_30_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_29 = qs_queue_29_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_28 = qs_queue_28_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_27 = qs_queue_27_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_26 = qs_queue_26_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_25 = qs_queue_25_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_24 = qs_queue_24_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_23 = qs_queue_23_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_22 = qs_queue_22_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_21 = qs_queue_21_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_20 = qs_queue_20_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_19 = qs_queue_19_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_18 = qs_queue_18_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_17 = qs_queue_17_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_16 = qs_queue_16_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_15 = qs_queue_15_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_14 = qs_queue_14_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_13 = qs_queue_13_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_12 = qs_queue_12_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_11 = qs_queue_11_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_10 = qs_queue_10_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_9 = qs_queue_9_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_8 = qs_queue_8_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_7 = qs_queue_7_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_6 = qs_queue_6_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_5 = qs_queue_5_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_4 = qs_queue_4_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_3 = qs_queue_3_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_2 = qs_queue_2_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_1 = qs_queue_1_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  enq_readys_0 = qs_queue_0_io_enq_ready; // @[Deinterleaver.scala 125:{33,33}]
  wire  _GEN_225 = 6'h1 == auto_out_rid ? enq_readys_1 : enq_readys_0; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_226 = 6'h2 == auto_out_rid ? enq_readys_2 : _GEN_225; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_227 = 6'h3 == auto_out_rid ? enq_readys_3 : _GEN_226; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_228 = 6'h4 == auto_out_rid ? enq_readys_4 : _GEN_227; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_229 = 6'h5 == auto_out_rid ? enq_readys_5 : _GEN_228; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_230 = 6'h6 == auto_out_rid ? enq_readys_6 : _GEN_229; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_231 = 6'h7 == auto_out_rid ? enq_readys_7 : _GEN_230; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_232 = 6'h8 == auto_out_rid ? enq_readys_8 : _GEN_231; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_233 = 6'h9 == auto_out_rid ? enq_readys_9 : _GEN_232; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_234 = 6'ha == auto_out_rid ? enq_readys_10 : _GEN_233; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_235 = 6'hb == auto_out_rid ? enq_readys_11 : _GEN_234; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_236 = 6'hc == auto_out_rid ? enq_readys_12 : _GEN_235; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_237 = 6'hd == auto_out_rid ? enq_readys_13 : _GEN_236; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_238 = 6'he == auto_out_rid ? enq_readys_14 : _GEN_237; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_239 = 6'hf == auto_out_rid ? enq_readys_15 : _GEN_238; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_240 = 6'h10 == auto_out_rid ? enq_readys_16 : _GEN_239; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_241 = 6'h11 == auto_out_rid ? enq_readys_17 : _GEN_240; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_242 = 6'h12 == auto_out_rid ? enq_readys_18 : _GEN_241; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_243 = 6'h13 == auto_out_rid ? enq_readys_19 : _GEN_242; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_244 = 6'h14 == auto_out_rid ? enq_readys_20 : _GEN_243; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_245 = 6'h15 == auto_out_rid ? enq_readys_21 : _GEN_244; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_246 = 6'h16 == auto_out_rid ? enq_readys_22 : _GEN_245; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_247 = 6'h17 == auto_out_rid ? enq_readys_23 : _GEN_246; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_248 = 6'h18 == auto_out_rid ? enq_readys_24 : _GEN_247; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_249 = 6'h19 == auto_out_rid ? enq_readys_25 : _GEN_248; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_250 = 6'h1a == auto_out_rid ? enq_readys_26 : _GEN_249; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_251 = 6'h1b == auto_out_rid ? enq_readys_27 : _GEN_250; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_252 = 6'h1c == auto_out_rid ? enq_readys_28 : _GEN_251; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_253 = 6'h1d == auto_out_rid ? enq_readys_29 : _GEN_252; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_254 = 6'h1e == auto_out_rid ? enq_readys_30 : _GEN_253; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_255 = 6'h1f == auto_out_rid ? enq_readys_31 : _GEN_254; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_256 = 6'h20 == auto_out_rid ? enq_readys_32 : _GEN_255; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_257 = 6'h21 == auto_out_rid ? enq_readys_33 : _GEN_256; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_258 = 6'h22 == auto_out_rid ? enq_readys_34 : _GEN_257; // @[Deinterleaver.scala 126:{21,21}]
  wire  _GEN_259 = 6'h23 == auto_out_rid ? enq_readys_35 : _GEN_258; // @[Deinterleaver.scala 126:{21,21}]
  wire  bundleOut_0_rready = 6'h24 == auto_out_rid ? enq_readys_36 : _GEN_259; // @[Deinterleaver.scala 126:{21,21}]
  wire  _pending_inc_T_1 = bundleOut_0_rready & auto_out_rvalid; // @[Decoupled.scala 50:35]
  wire  pending_inc = enq_OH[0] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  _pending_dec_T_1 = auto_in_rready & locked; // @[Decoupled.scala 50:35]
  wire  deq_bits_36_last = qs_queue_36_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_35_last = qs_queue_35_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_34_last = qs_queue_34_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_33_last = qs_queue_33_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_32_last = qs_queue_32_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_31_last = qs_queue_31_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_30_last = qs_queue_30_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_29_last = qs_queue_29_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_28_last = qs_queue_28_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_27_last = qs_queue_27_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_26_last = qs_queue_26_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_25_last = qs_queue_25_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_24_last = qs_queue_24_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_23_last = qs_queue_23_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_22_last = qs_queue_22_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_21_last = qs_queue_21_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_20_last = qs_queue_20_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_19_last = qs_queue_19_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_18_last = qs_queue_18_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_17_last = qs_queue_17_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_16_last = qs_queue_16_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_15_last = qs_queue_15_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_14_last = qs_queue_14_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_13_last = qs_queue_13_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_12_last = qs_queue_12_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_11_last = qs_queue_11_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_10_last = qs_queue_10_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_9_last = qs_queue_9_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_8_last = qs_queue_8_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_7_last = qs_queue_7_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_6_last = qs_queue_6_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_5_last = qs_queue_5_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_4_last = qs_queue_4_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_3_last = qs_queue_3_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_2_last = qs_queue_2_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_1_last = qs_queue_1_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  deq_bits_0_last = qs_queue_0_io_deq_bits_last; // @[Deinterleaver.scala 114:{31,31}]
  wire  _GEN_3 = 6'h1 == deq_id ? deq_bits_1_last : deq_bits_0_last; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_4 = 6'h2 == deq_id ? deq_bits_2_last : _GEN_3; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_5 = 6'h3 == deq_id ? deq_bits_3_last : _GEN_4; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_6 = 6'h4 == deq_id ? deq_bits_4_last : _GEN_5; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_7 = 6'h5 == deq_id ? deq_bits_5_last : _GEN_6; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_8 = 6'h6 == deq_id ? deq_bits_6_last : _GEN_7; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_9 = 6'h7 == deq_id ? deq_bits_7_last : _GEN_8; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_10 = 6'h8 == deq_id ? deq_bits_8_last : _GEN_9; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_11 = 6'h9 == deq_id ? deq_bits_9_last : _GEN_10; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_12 = 6'ha == deq_id ? deq_bits_10_last : _GEN_11; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_13 = 6'hb == deq_id ? deq_bits_11_last : _GEN_12; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_14 = 6'hc == deq_id ? deq_bits_12_last : _GEN_13; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_15 = 6'hd == deq_id ? deq_bits_13_last : _GEN_14; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_16 = 6'he == deq_id ? deq_bits_14_last : _GEN_15; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_17 = 6'hf == deq_id ? deq_bits_15_last : _GEN_16; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_18 = 6'h10 == deq_id ? deq_bits_16_last : _GEN_17; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_19 = 6'h11 == deq_id ? deq_bits_17_last : _GEN_18; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_20 = 6'h12 == deq_id ? deq_bits_18_last : _GEN_19; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_21 = 6'h13 == deq_id ? deq_bits_19_last : _GEN_20; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_22 = 6'h14 == deq_id ? deq_bits_20_last : _GEN_21; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_23 = 6'h15 == deq_id ? deq_bits_21_last : _GEN_22; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_24 = 6'h16 == deq_id ? deq_bits_22_last : _GEN_23; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_25 = 6'h17 == deq_id ? deq_bits_23_last : _GEN_24; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_26 = 6'h18 == deq_id ? deq_bits_24_last : _GEN_25; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_27 = 6'h19 == deq_id ? deq_bits_25_last : _GEN_26; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_28 = 6'h1a == deq_id ? deq_bits_26_last : _GEN_27; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_29 = 6'h1b == deq_id ? deq_bits_27_last : _GEN_28; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_30 = 6'h1c == deq_id ? deq_bits_28_last : _GEN_29; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_31 = 6'h1d == deq_id ? deq_bits_29_last : _GEN_30; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_32 = 6'h1e == deq_id ? deq_bits_30_last : _GEN_31; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_33 = 6'h1f == deq_id ? deq_bits_31_last : _GEN_32; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_34 = 6'h20 == deq_id ? deq_bits_32_last : _GEN_33; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_35 = 6'h21 == deq_id ? deq_bits_33_last : _GEN_34; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_36 = 6'h22 == deq_id ? deq_bits_34_last : _GEN_35; // @[Deinterleaver.scala 115:{20,20}]
  wire  _GEN_37 = 6'h23 == deq_id ? deq_bits_35_last : _GEN_36; // @[Deinterleaver.scala 115:{20,20}]
  wire  bundleIn_0_rlast = 6'h24 == deq_id ? deq_bits_36_last : _GEN_37; // @[Deinterleaver.scala 115:{20,20}]
  wire  pending_dec = deq_OH[0] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_261 = {{1'd0}, pending_inc}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_1 = pending_count + _GEN_261; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_262 = {{1'd0}, pending_dec}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next = _pending_next_T_1 - _GEN_262; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_12 = pending_next != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_1; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_1 = enq_OH[1] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_1 = deq_OH[1] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_263 = {{1'd0}, pending_inc_1}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_5 = pending_count_1 + _GEN_263; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_264 = {{1'd0}, pending_dec_1}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_1 = _pending_next_T_5 - _GEN_264; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_25 = pending_next_1 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_2; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_2 = enq_OH[2] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_2 = deq_OH[2] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_265 = {{1'd0}, pending_inc_2}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_9 = pending_count_2 + _GEN_265; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_266 = {{1'd0}, pending_dec_2}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_2 = _pending_next_T_9 - _GEN_266; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_38 = pending_next_2 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_3; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_3 = enq_OH[3] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_3 = deq_OH[3] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_267 = {{1'd0}, pending_inc_3}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_13 = pending_count_3 + _GEN_267; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_268 = {{1'd0}, pending_dec_3}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_3 = _pending_next_T_13 - _GEN_268; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_51 = pending_next_3 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_4; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_4 = enq_OH[4] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_4 = deq_OH[4] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_269 = {{1'd0}, pending_inc_4}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_17 = pending_count_4 + _GEN_269; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_270 = {{1'd0}, pending_dec_4}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_4 = _pending_next_T_17 - _GEN_270; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_64 = pending_next_4 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_5; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_5 = enq_OH[5] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_5 = deq_OH[5] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_271 = {{1'd0}, pending_inc_5}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_21 = pending_count_5 + _GEN_271; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_272 = {{1'd0}, pending_dec_5}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_5 = _pending_next_T_21 - _GEN_272; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_77 = pending_next_5 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_6; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_6 = enq_OH[6] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_6 = deq_OH[6] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_273 = {{1'd0}, pending_inc_6}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_25 = pending_count_6 + _GEN_273; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_274 = {{1'd0}, pending_dec_6}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_6 = _pending_next_T_25 - _GEN_274; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_90 = pending_next_6 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_7; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_7 = enq_OH[7] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_7 = deq_OH[7] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_275 = {{1'd0}, pending_inc_7}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_29 = pending_count_7 + _GEN_275; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_276 = {{1'd0}, pending_dec_7}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_7 = _pending_next_T_29 - _GEN_276; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_103 = pending_next_7 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_8; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_8 = enq_OH[8] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_8 = deq_OH[8] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_277 = {{1'd0}, pending_inc_8}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_33 = pending_count_8 + _GEN_277; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_278 = {{1'd0}, pending_dec_8}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_8 = _pending_next_T_33 - _GEN_278; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_116 = pending_next_8 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_9; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_9 = enq_OH[9] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_9 = deq_OH[9] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_279 = {{1'd0}, pending_inc_9}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_37 = pending_count_9 + _GEN_279; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_280 = {{1'd0}, pending_dec_9}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_9 = _pending_next_T_37 - _GEN_280; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_129 = pending_next_9 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_10; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_10 = enq_OH[10] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_10 = deq_OH[10] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_281 = {{1'd0}, pending_inc_10}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_41 = pending_count_10 + _GEN_281; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_282 = {{1'd0}, pending_dec_10}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_10 = _pending_next_T_41 - _GEN_282; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_142 = pending_next_10 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_11; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_11 = enq_OH[11] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_11 = deq_OH[11] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_283 = {{1'd0}, pending_inc_11}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_45 = pending_count_11 + _GEN_283; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_284 = {{1'd0}, pending_dec_11}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_11 = _pending_next_T_45 - _GEN_284; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_155 = pending_next_11 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_12; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_12 = enq_OH[12] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_12 = deq_OH[12] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_285 = {{1'd0}, pending_inc_12}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_49 = pending_count_12 + _GEN_285; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_286 = {{1'd0}, pending_dec_12}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_12 = _pending_next_T_49 - _GEN_286; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_168 = pending_next_12 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_13; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_13 = enq_OH[13] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_13 = deq_OH[13] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_287 = {{1'd0}, pending_inc_13}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_53 = pending_count_13 + _GEN_287; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_288 = {{1'd0}, pending_dec_13}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_13 = _pending_next_T_53 - _GEN_288; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_181 = pending_next_13 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_14; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_14 = enq_OH[14] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_14 = deq_OH[14] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_289 = {{1'd0}, pending_inc_14}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_57 = pending_count_14 + _GEN_289; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_290 = {{1'd0}, pending_dec_14}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_14 = _pending_next_T_57 - _GEN_290; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_194 = pending_next_14 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_15; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_15 = enq_OH[15] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_15 = deq_OH[15] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_291 = {{1'd0}, pending_inc_15}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_61 = pending_count_15 + _GEN_291; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_292 = {{1'd0}, pending_dec_15}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_15 = _pending_next_T_61 - _GEN_292; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_207 = pending_next_15 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_16; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_16 = enq_OH[16] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_16 = deq_OH[16] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_293 = {{1'd0}, pending_inc_16}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_65 = pending_count_16 + _GEN_293; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_294 = {{1'd0}, pending_dec_16}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_16 = _pending_next_T_65 - _GEN_294; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_220 = pending_next_16 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_17; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_17 = enq_OH[17] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_17 = deq_OH[17] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_295 = {{1'd0}, pending_inc_17}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_69 = pending_count_17 + _GEN_295; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_296 = {{1'd0}, pending_dec_17}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_17 = _pending_next_T_69 - _GEN_296; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_233 = pending_next_17 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_18; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_18 = enq_OH[18] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_18 = deq_OH[18] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_297 = {{1'd0}, pending_inc_18}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_73 = pending_count_18 + _GEN_297; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_298 = {{1'd0}, pending_dec_18}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_18 = _pending_next_T_73 - _GEN_298; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_246 = pending_next_18 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_19; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_19 = enq_OH[19] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_19 = deq_OH[19] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_299 = {{1'd0}, pending_inc_19}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_77 = pending_count_19 + _GEN_299; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_300 = {{1'd0}, pending_dec_19}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_19 = _pending_next_T_77 - _GEN_300; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_259 = pending_next_19 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_20; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_20 = enq_OH[20] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_20 = deq_OH[20] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_301 = {{1'd0}, pending_inc_20}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_81 = pending_count_20 + _GEN_301; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_302 = {{1'd0}, pending_dec_20}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_20 = _pending_next_T_81 - _GEN_302; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_272 = pending_next_20 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_21; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_21 = enq_OH[21] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_21 = deq_OH[21] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_303 = {{1'd0}, pending_inc_21}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_85 = pending_count_21 + _GEN_303; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_304 = {{1'd0}, pending_dec_21}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_21 = _pending_next_T_85 - _GEN_304; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_285 = pending_next_21 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_22; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_22 = enq_OH[22] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_22 = deq_OH[22] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_305 = {{1'd0}, pending_inc_22}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_89 = pending_count_22 + _GEN_305; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_306 = {{1'd0}, pending_dec_22}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_22 = _pending_next_T_89 - _GEN_306; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_298 = pending_next_22 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_23; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_23 = enq_OH[23] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_23 = deq_OH[23] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_307 = {{1'd0}, pending_inc_23}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_93 = pending_count_23 + _GEN_307; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_308 = {{1'd0}, pending_dec_23}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_23 = _pending_next_T_93 - _GEN_308; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_311 = pending_next_23 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_24; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_24 = enq_OH[24] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_24 = deq_OH[24] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_309 = {{1'd0}, pending_inc_24}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_97 = pending_count_24 + _GEN_309; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_310 = {{1'd0}, pending_dec_24}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_24 = _pending_next_T_97 - _GEN_310; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_324 = pending_next_24 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_25; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_25 = enq_OH[25] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_25 = deq_OH[25] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_311 = {{1'd0}, pending_inc_25}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_101 = pending_count_25 + _GEN_311; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_312 = {{1'd0}, pending_dec_25}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_25 = _pending_next_T_101 - _GEN_312; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_337 = pending_next_25 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_26; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_26 = enq_OH[26] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_26 = deq_OH[26] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_313 = {{1'd0}, pending_inc_26}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_105 = pending_count_26 + _GEN_313; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_314 = {{1'd0}, pending_dec_26}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_26 = _pending_next_T_105 - _GEN_314; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_350 = pending_next_26 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_27; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_27 = enq_OH[27] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_27 = deq_OH[27] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_315 = {{1'd0}, pending_inc_27}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_109 = pending_count_27 + _GEN_315; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_316 = {{1'd0}, pending_dec_27}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_27 = _pending_next_T_109 - _GEN_316; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_363 = pending_next_27 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_28; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_28 = enq_OH[28] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_28 = deq_OH[28] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_317 = {{1'd0}, pending_inc_28}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_113 = pending_count_28 + _GEN_317; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_318 = {{1'd0}, pending_dec_28}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_28 = _pending_next_T_113 - _GEN_318; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_376 = pending_next_28 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_29; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_29 = enq_OH[29] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_29 = deq_OH[29] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_319 = {{1'd0}, pending_inc_29}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_117 = pending_count_29 + _GEN_319; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_320 = {{1'd0}, pending_dec_29}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_29 = _pending_next_T_117 - _GEN_320; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_389 = pending_next_29 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_30; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_30 = enq_OH[30] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_30 = deq_OH[30] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_321 = {{1'd0}, pending_inc_30}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_121 = pending_count_30 + _GEN_321; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_322 = {{1'd0}, pending_dec_30}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_30 = _pending_next_T_121 - _GEN_322; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_402 = pending_next_30 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_31; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_31 = enq_OH[31] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_31 = deq_OH[31] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_323 = {{1'd0}, pending_inc_31}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_125 = pending_count_31 + _GEN_323; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_324 = {{1'd0}, pending_dec_31}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_31 = _pending_next_T_125 - _GEN_324; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_415 = pending_next_31 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_32; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_32 = enq_OH[32] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_32 = deq_OH[32] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_325 = {{1'd0}, pending_inc_32}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_129 = pending_count_32 + _GEN_325; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_326 = {{1'd0}, pending_dec_32}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_32 = _pending_next_T_129 - _GEN_326; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_428 = pending_next_32 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_33; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_33 = enq_OH[33] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_33 = deq_OH[33] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_327 = {{1'd0}, pending_inc_33}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_133 = pending_count_33 + _GEN_327; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_328 = {{1'd0}, pending_dec_33}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_33 = _pending_next_T_133 - _GEN_328; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_441 = pending_next_33 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_34; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_34 = enq_OH[34] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_34 = deq_OH[34] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_329 = {{1'd0}, pending_inc_34}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_137 = pending_count_34 + _GEN_329; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_330 = {{1'd0}, pending_dec_34}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_34 = _pending_next_T_137 - _GEN_330; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_454 = pending_next_34 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_35; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_35 = enq_OH[35] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_35 = deq_OH[35] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_331 = {{1'd0}, pending_inc_35}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_141 = pending_count_35 + _GEN_331; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_332 = {{1'd0}, pending_dec_35}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_35 = _pending_next_T_141 - _GEN_332; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_467 = pending_next_35 != 2'h0; // @[Deinterleaver.scala 101:18]
  reg [1:0] pending_count_36; // @[Deinterleaver.scala 92:32]
  wire  pending_inc_36 = enq_OH[36] & _pending_inc_T_1 & auto_out_rlast; // @[Deinterleaver.scala 94:49]
  wire  pending_dec_36 = deq_OH[36] & _pending_dec_T_1 & bundleIn_0_rlast; // @[Deinterleaver.scala 95:48]
  wire [1:0] _GEN_333 = {{1'd0}, pending_inc_36}; // @[Deinterleaver.scala 96:27]
  wire [1:0] _pending_next_T_145 = pending_count_36 + _GEN_333; // @[Deinterleaver.scala 96:27]
  wire [1:0] _GEN_334 = {{1'd0}, pending_dec_36}; // @[Deinterleaver.scala 96:40]
  wire [1:0] pending_next_36 = _pending_next_T_145 - _GEN_334; // @[Deinterleaver.scala 96:40]
  wire  _pending_T_480 = pending_next_36 != 2'h0; // @[Deinterleaver.scala 101:18]
  wire [8:0] pending_lo_lo = {_pending_T_116,_pending_T_103,_pending_T_90,_pending_T_77,_pending_T_64,_pending_T_51,
    _pending_T_38,_pending_T_25,_pending_T_12}; // @[Cat.scala 31:58]
  wire [17:0] pending_lo = {_pending_T_233,_pending_T_220,_pending_T_207,_pending_T_194,_pending_T_181,_pending_T_168,
    _pending_T_155,_pending_T_142,_pending_T_129,pending_lo_lo}; // @[Cat.scala 31:58]
  wire [9:0] pending_hi_hi = {_pending_T_480,_pending_T_467,_pending_T_454,_pending_T_441,_pending_T_428,_pending_T_415,
    _pending_T_402,_pending_T_389,_pending_T_376,_pending_T_363}; // @[Cat.scala 31:58]
  wire [18:0] pending_hi = {pending_hi_hi,_pending_T_350,_pending_T_337,_pending_T_324,_pending_T_311,_pending_T_298,
    _pending_T_285,_pending_T_272,_pending_T_259,_pending_T_246}; // @[Cat.scala 31:58]
  wire [36:0] pending = {pending_hi,pending_lo}; // @[Cat.scala 31:58]
  wire [37:0] _winner_T = {pending, 1'h0}; // @[package.scala 244:48]
  wire [36:0] _winner_T_2 = pending | _winner_T[36:0]; // @[package.scala 244:43]
  wire [38:0] _winner_T_3 = {_winner_T_2, 2'h0}; // @[package.scala 244:48]
  wire [36:0] _winner_T_5 = _winner_T_2 | _winner_T_3[36:0]; // @[package.scala 244:43]
  wire [40:0] _winner_T_6 = {_winner_T_5, 4'h0}; // @[package.scala 244:48]
  wire [36:0] _winner_T_8 = _winner_T_5 | _winner_T_6[36:0]; // @[package.scala 244:43]
  wire [44:0] _winner_T_9 = {_winner_T_8, 8'h0}; // @[package.scala 244:48]
  wire [36:0] _winner_T_11 = _winner_T_8 | _winner_T_9[36:0]; // @[package.scala 244:43]
  wire [52:0] _winner_T_12 = {_winner_T_11, 16'h0}; // @[package.scala 244:48]
  wire [36:0] _winner_T_14 = _winner_T_11 | _winner_T_12[36:0]; // @[package.scala 244:43]
  wire [68:0] _winner_T_15 = {_winner_T_14, 32'h0}; // @[package.scala 244:48]
  wire [36:0] _winner_T_17 = _winner_T_14 | _winner_T_15[36:0]; // @[package.scala 244:43]
  wire [37:0] _winner_T_19 = {_winner_T_17, 1'h0}; // @[Deinterleaver.scala 106:51]
  wire [37:0] _winner_T_20 = ~_winner_T_19; // @[Deinterleaver.scala 106:33]
  wire [37:0] _GEN_335 = {{1'd0}, pending}; // @[Deinterleaver.scala 106:31]
  wire [37:0] winner = _GEN_335 & _winner_T_20; // @[Deinterleaver.scala 106:31]
  wire [5:0] deq_id_hi = winner[37:32]; // @[OneHot.scala 30:18]
  wire [31:0] deq_id_lo = winner[31:0]; // @[OneHot.scala 31:18]
  wire  _deq_id_T = |deq_id_hi; // @[OneHot.scala 32:14]
  wire [31:0] _GEN_336 = {{26'd0}, deq_id_hi}; // @[OneHot.scala 32:28]
  wire [31:0] _deq_id_T_1 = _GEN_336 | deq_id_lo; // @[OneHot.scala 32:28]
  wire [15:0] deq_id_hi_1 = _deq_id_T_1[31:16]; // @[OneHot.scala 30:18]
  wire [15:0] deq_id_lo_1 = _deq_id_T_1[15:0]; // @[OneHot.scala 31:18]
  wire  _deq_id_T_2 = |deq_id_hi_1; // @[OneHot.scala 32:14]
  wire [15:0] _deq_id_T_3 = deq_id_hi_1 | deq_id_lo_1; // @[OneHot.scala 32:28]
  wire [7:0] deq_id_hi_2 = _deq_id_T_3[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] deq_id_lo_2 = _deq_id_T_3[7:0]; // @[OneHot.scala 31:18]
  wire  _deq_id_T_4 = |deq_id_hi_2; // @[OneHot.scala 32:14]
  wire [7:0] _deq_id_T_5 = deq_id_hi_2 | deq_id_lo_2; // @[OneHot.scala 32:28]
  wire [3:0] deq_id_hi_3 = _deq_id_T_5[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] deq_id_lo_3 = _deq_id_T_5[3:0]; // @[OneHot.scala 31:18]
  wire  _deq_id_T_6 = |deq_id_hi_3; // @[OneHot.scala 32:14]
  wire [3:0] _deq_id_T_7 = deq_id_hi_3 | deq_id_lo_3; // @[OneHot.scala 32:28]
  wire [1:0] deq_id_hi_4 = _deq_id_T_7[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] deq_id_lo_4 = _deq_id_T_7[1:0]; // @[OneHot.scala 31:18]
  wire  _deq_id_T_8 = |deq_id_hi_4; // @[OneHot.scala 32:14]
  wire [1:0] _deq_id_T_9 = deq_id_hi_4 | deq_id_lo_4; // @[OneHot.scala 32:28]
  wire [5:0] _deq_id_T_15 = {_deq_id_T,_deq_id_T_2,_deq_id_T_4,_deq_id_T_6,_deq_id_T_8,_deq_id_T_9[1]}; // @[Cat.scala 31:58]
  wire [5:0] deq_bits_0_echo_tl_state_source = qs_queue_0_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] deq_bits_1_echo_tl_state_source = qs_queue_1_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_40 = 6'h1 == deq_id ? deq_bits_1_echo_tl_state_source : deq_bits_0_echo_tl_state_source; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_2_echo_tl_state_source = qs_queue_2_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_41 = 6'h2 == deq_id ? deq_bits_2_echo_tl_state_source : _GEN_40; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_3_echo_tl_state_source = qs_queue_3_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_42 = 6'h3 == deq_id ? deq_bits_3_echo_tl_state_source : _GEN_41; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_4_echo_tl_state_source = qs_queue_4_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_43 = 6'h4 == deq_id ? deq_bits_4_echo_tl_state_source : _GEN_42; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_5_echo_tl_state_source = qs_queue_5_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_44 = 6'h5 == deq_id ? deq_bits_5_echo_tl_state_source : _GEN_43; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_6_echo_tl_state_source = qs_queue_6_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_45 = 6'h6 == deq_id ? deq_bits_6_echo_tl_state_source : _GEN_44; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_7_echo_tl_state_source = qs_queue_7_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_46 = 6'h7 == deq_id ? deq_bits_7_echo_tl_state_source : _GEN_45; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_8_echo_tl_state_source = qs_queue_8_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_47 = 6'h8 == deq_id ? deq_bits_8_echo_tl_state_source : _GEN_46; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_9_echo_tl_state_source = qs_queue_9_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_48 = 6'h9 == deq_id ? deq_bits_9_echo_tl_state_source : _GEN_47; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_10_echo_tl_state_source = qs_queue_10_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_49 = 6'ha == deq_id ? deq_bits_10_echo_tl_state_source : _GEN_48; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_11_echo_tl_state_source = qs_queue_11_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_50 = 6'hb == deq_id ? deq_bits_11_echo_tl_state_source : _GEN_49; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_12_echo_tl_state_source = qs_queue_12_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_51 = 6'hc == deq_id ? deq_bits_12_echo_tl_state_source : _GEN_50; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_13_echo_tl_state_source = qs_queue_13_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_52 = 6'hd == deq_id ? deq_bits_13_echo_tl_state_source : _GEN_51; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_14_echo_tl_state_source = qs_queue_14_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_53 = 6'he == deq_id ? deq_bits_14_echo_tl_state_source : _GEN_52; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_15_echo_tl_state_source = qs_queue_15_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_54 = 6'hf == deq_id ? deq_bits_15_echo_tl_state_source : _GEN_53; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_16_echo_tl_state_source = qs_queue_16_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_55 = 6'h10 == deq_id ? deq_bits_16_echo_tl_state_source : _GEN_54; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_17_echo_tl_state_source = qs_queue_17_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_56 = 6'h11 == deq_id ? deq_bits_17_echo_tl_state_source : _GEN_55; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_18_echo_tl_state_source = qs_queue_18_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_57 = 6'h12 == deq_id ? deq_bits_18_echo_tl_state_source : _GEN_56; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_19_echo_tl_state_source = qs_queue_19_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_58 = 6'h13 == deq_id ? deq_bits_19_echo_tl_state_source : _GEN_57; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_20_echo_tl_state_source = qs_queue_20_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_59 = 6'h14 == deq_id ? deq_bits_20_echo_tl_state_source : _GEN_58; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_21_echo_tl_state_source = qs_queue_21_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_60 = 6'h15 == deq_id ? deq_bits_21_echo_tl_state_source : _GEN_59; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_22_echo_tl_state_source = qs_queue_22_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_61 = 6'h16 == deq_id ? deq_bits_22_echo_tl_state_source : _GEN_60; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_23_echo_tl_state_source = qs_queue_23_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_62 = 6'h17 == deq_id ? deq_bits_23_echo_tl_state_source : _GEN_61; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_24_echo_tl_state_source = qs_queue_24_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_63 = 6'h18 == deq_id ? deq_bits_24_echo_tl_state_source : _GEN_62; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_25_echo_tl_state_source = qs_queue_25_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_64 = 6'h19 == deq_id ? deq_bits_25_echo_tl_state_source : _GEN_63; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_26_echo_tl_state_source = qs_queue_26_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_65 = 6'h1a == deq_id ? deq_bits_26_echo_tl_state_source : _GEN_64; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_27_echo_tl_state_source = qs_queue_27_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_66 = 6'h1b == deq_id ? deq_bits_27_echo_tl_state_source : _GEN_65; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_28_echo_tl_state_source = qs_queue_28_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_67 = 6'h1c == deq_id ? deq_bits_28_echo_tl_state_source : _GEN_66; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_29_echo_tl_state_source = qs_queue_29_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_68 = 6'h1d == deq_id ? deq_bits_29_echo_tl_state_source : _GEN_67; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_30_echo_tl_state_source = qs_queue_30_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_69 = 6'h1e == deq_id ? deq_bits_30_echo_tl_state_source : _GEN_68; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_31_echo_tl_state_source = qs_queue_31_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_70 = 6'h1f == deq_id ? deq_bits_31_echo_tl_state_source : _GEN_69; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_32_echo_tl_state_source = qs_queue_32_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_71 = 6'h20 == deq_id ? deq_bits_32_echo_tl_state_source : _GEN_70; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_33_echo_tl_state_source = qs_queue_33_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_72 = 6'h21 == deq_id ? deq_bits_33_echo_tl_state_source : _GEN_71; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_34_echo_tl_state_source = qs_queue_34_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_73 = 6'h22 == deq_id ? deq_bits_34_echo_tl_state_source : _GEN_72; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_35_echo_tl_state_source = qs_queue_35_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_74 = 6'h23 == deq_id ? deq_bits_35_echo_tl_state_source : _GEN_73; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_36_echo_tl_state_source = qs_queue_36_io_deq_bits_echo_tl_state_source; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] deq_bits_0_echo_tl_state_size = qs_queue_0_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] deq_bits_1_echo_tl_state_size = qs_queue_1_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_77 = 6'h1 == deq_id ? deq_bits_1_echo_tl_state_size : deq_bits_0_echo_tl_state_size; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_2_echo_tl_state_size = qs_queue_2_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_78 = 6'h2 == deq_id ? deq_bits_2_echo_tl_state_size : _GEN_77; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_3_echo_tl_state_size = qs_queue_3_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_79 = 6'h3 == deq_id ? deq_bits_3_echo_tl_state_size : _GEN_78; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_4_echo_tl_state_size = qs_queue_4_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_80 = 6'h4 == deq_id ? deq_bits_4_echo_tl_state_size : _GEN_79; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_5_echo_tl_state_size = qs_queue_5_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_81 = 6'h5 == deq_id ? deq_bits_5_echo_tl_state_size : _GEN_80; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_6_echo_tl_state_size = qs_queue_6_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_82 = 6'h6 == deq_id ? deq_bits_6_echo_tl_state_size : _GEN_81; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_7_echo_tl_state_size = qs_queue_7_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_83 = 6'h7 == deq_id ? deq_bits_7_echo_tl_state_size : _GEN_82; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_8_echo_tl_state_size = qs_queue_8_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_84 = 6'h8 == deq_id ? deq_bits_8_echo_tl_state_size : _GEN_83; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_9_echo_tl_state_size = qs_queue_9_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_85 = 6'h9 == deq_id ? deq_bits_9_echo_tl_state_size : _GEN_84; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_10_echo_tl_state_size = qs_queue_10_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_86 = 6'ha == deq_id ? deq_bits_10_echo_tl_state_size : _GEN_85; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_11_echo_tl_state_size = qs_queue_11_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_87 = 6'hb == deq_id ? deq_bits_11_echo_tl_state_size : _GEN_86; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_12_echo_tl_state_size = qs_queue_12_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_88 = 6'hc == deq_id ? deq_bits_12_echo_tl_state_size : _GEN_87; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_13_echo_tl_state_size = qs_queue_13_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_89 = 6'hd == deq_id ? deq_bits_13_echo_tl_state_size : _GEN_88; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_14_echo_tl_state_size = qs_queue_14_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_90 = 6'he == deq_id ? deq_bits_14_echo_tl_state_size : _GEN_89; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_15_echo_tl_state_size = qs_queue_15_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_91 = 6'hf == deq_id ? deq_bits_15_echo_tl_state_size : _GEN_90; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_16_echo_tl_state_size = qs_queue_16_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_92 = 6'h10 == deq_id ? deq_bits_16_echo_tl_state_size : _GEN_91; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_17_echo_tl_state_size = qs_queue_17_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_93 = 6'h11 == deq_id ? deq_bits_17_echo_tl_state_size : _GEN_92; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_18_echo_tl_state_size = qs_queue_18_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_94 = 6'h12 == deq_id ? deq_bits_18_echo_tl_state_size : _GEN_93; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_19_echo_tl_state_size = qs_queue_19_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_95 = 6'h13 == deq_id ? deq_bits_19_echo_tl_state_size : _GEN_94; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_20_echo_tl_state_size = qs_queue_20_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_96 = 6'h14 == deq_id ? deq_bits_20_echo_tl_state_size : _GEN_95; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_21_echo_tl_state_size = qs_queue_21_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_97 = 6'h15 == deq_id ? deq_bits_21_echo_tl_state_size : _GEN_96; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_22_echo_tl_state_size = qs_queue_22_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_98 = 6'h16 == deq_id ? deq_bits_22_echo_tl_state_size : _GEN_97; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_23_echo_tl_state_size = qs_queue_23_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_99 = 6'h17 == deq_id ? deq_bits_23_echo_tl_state_size : _GEN_98; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_24_echo_tl_state_size = qs_queue_24_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_100 = 6'h18 == deq_id ? deq_bits_24_echo_tl_state_size : _GEN_99; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_25_echo_tl_state_size = qs_queue_25_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_101 = 6'h19 == deq_id ? deq_bits_25_echo_tl_state_size : _GEN_100; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_26_echo_tl_state_size = qs_queue_26_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_102 = 6'h1a == deq_id ? deq_bits_26_echo_tl_state_size : _GEN_101; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_27_echo_tl_state_size = qs_queue_27_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_103 = 6'h1b == deq_id ? deq_bits_27_echo_tl_state_size : _GEN_102; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_28_echo_tl_state_size = qs_queue_28_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_104 = 6'h1c == deq_id ? deq_bits_28_echo_tl_state_size : _GEN_103; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_29_echo_tl_state_size = qs_queue_29_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_105 = 6'h1d == deq_id ? deq_bits_29_echo_tl_state_size : _GEN_104; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_30_echo_tl_state_size = qs_queue_30_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_106 = 6'h1e == deq_id ? deq_bits_30_echo_tl_state_size : _GEN_105; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_31_echo_tl_state_size = qs_queue_31_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_107 = 6'h1f == deq_id ? deq_bits_31_echo_tl_state_size : _GEN_106; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_32_echo_tl_state_size = qs_queue_32_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_108 = 6'h20 == deq_id ? deq_bits_32_echo_tl_state_size : _GEN_107; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_33_echo_tl_state_size = qs_queue_33_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_109 = 6'h21 == deq_id ? deq_bits_33_echo_tl_state_size : _GEN_108; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_34_echo_tl_state_size = qs_queue_34_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_110 = 6'h22 == deq_id ? deq_bits_34_echo_tl_state_size : _GEN_109; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_35_echo_tl_state_size = qs_queue_35_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [3:0] _GEN_111 = 6'h23 == deq_id ? deq_bits_35_echo_tl_state_size : _GEN_110; // @[Deinterleaver.scala 115:{20,20}]
  wire [3:0] deq_bits_36_echo_tl_state_size = qs_queue_36_io_deq_bits_echo_tl_state_size; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] deq_bits_0_resp = qs_queue_0_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] deq_bits_1_resp = qs_queue_1_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_114 = 6'h1 == deq_id ? deq_bits_1_resp : deq_bits_0_resp; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_2_resp = qs_queue_2_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_115 = 6'h2 == deq_id ? deq_bits_2_resp : _GEN_114; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_3_resp = qs_queue_3_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_116 = 6'h3 == deq_id ? deq_bits_3_resp : _GEN_115; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_4_resp = qs_queue_4_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_117 = 6'h4 == deq_id ? deq_bits_4_resp : _GEN_116; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_5_resp = qs_queue_5_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_118 = 6'h5 == deq_id ? deq_bits_5_resp : _GEN_117; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_6_resp = qs_queue_6_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_119 = 6'h6 == deq_id ? deq_bits_6_resp : _GEN_118; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_7_resp = qs_queue_7_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_120 = 6'h7 == deq_id ? deq_bits_7_resp : _GEN_119; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_8_resp = qs_queue_8_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_121 = 6'h8 == deq_id ? deq_bits_8_resp : _GEN_120; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_9_resp = qs_queue_9_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_122 = 6'h9 == deq_id ? deq_bits_9_resp : _GEN_121; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_10_resp = qs_queue_10_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_123 = 6'ha == deq_id ? deq_bits_10_resp : _GEN_122; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_11_resp = qs_queue_11_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_124 = 6'hb == deq_id ? deq_bits_11_resp : _GEN_123; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_12_resp = qs_queue_12_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_125 = 6'hc == deq_id ? deq_bits_12_resp : _GEN_124; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_13_resp = qs_queue_13_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_126 = 6'hd == deq_id ? deq_bits_13_resp : _GEN_125; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_14_resp = qs_queue_14_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_127 = 6'he == deq_id ? deq_bits_14_resp : _GEN_126; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_15_resp = qs_queue_15_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_128 = 6'hf == deq_id ? deq_bits_15_resp : _GEN_127; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_16_resp = qs_queue_16_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_129 = 6'h10 == deq_id ? deq_bits_16_resp : _GEN_128; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_17_resp = qs_queue_17_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_130 = 6'h11 == deq_id ? deq_bits_17_resp : _GEN_129; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_18_resp = qs_queue_18_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_131 = 6'h12 == deq_id ? deq_bits_18_resp : _GEN_130; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_19_resp = qs_queue_19_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_132 = 6'h13 == deq_id ? deq_bits_19_resp : _GEN_131; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_20_resp = qs_queue_20_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_133 = 6'h14 == deq_id ? deq_bits_20_resp : _GEN_132; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_21_resp = qs_queue_21_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_134 = 6'h15 == deq_id ? deq_bits_21_resp : _GEN_133; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_22_resp = qs_queue_22_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_135 = 6'h16 == deq_id ? deq_bits_22_resp : _GEN_134; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_23_resp = qs_queue_23_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_136 = 6'h17 == deq_id ? deq_bits_23_resp : _GEN_135; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_24_resp = qs_queue_24_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_137 = 6'h18 == deq_id ? deq_bits_24_resp : _GEN_136; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_25_resp = qs_queue_25_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_138 = 6'h19 == deq_id ? deq_bits_25_resp : _GEN_137; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_26_resp = qs_queue_26_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_139 = 6'h1a == deq_id ? deq_bits_26_resp : _GEN_138; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_27_resp = qs_queue_27_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_140 = 6'h1b == deq_id ? deq_bits_27_resp : _GEN_139; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_28_resp = qs_queue_28_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_141 = 6'h1c == deq_id ? deq_bits_28_resp : _GEN_140; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_29_resp = qs_queue_29_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_142 = 6'h1d == deq_id ? deq_bits_29_resp : _GEN_141; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_30_resp = qs_queue_30_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_143 = 6'h1e == deq_id ? deq_bits_30_resp : _GEN_142; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_31_resp = qs_queue_31_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_144 = 6'h1f == deq_id ? deq_bits_31_resp : _GEN_143; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_32_resp = qs_queue_32_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_145 = 6'h20 == deq_id ? deq_bits_32_resp : _GEN_144; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_33_resp = qs_queue_33_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_146 = 6'h21 == deq_id ? deq_bits_33_resp : _GEN_145; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_34_resp = qs_queue_34_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_147 = 6'h22 == deq_id ? deq_bits_34_resp : _GEN_146; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_35_resp = qs_queue_35_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [1:0] _GEN_148 = 6'h23 == deq_id ? deq_bits_35_resp : _GEN_147; // @[Deinterleaver.scala 115:{20,20}]
  wire [1:0] deq_bits_36_resp = qs_queue_36_io_deq_bits_resp; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] deq_bits_0_data = qs_queue_0_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] deq_bits_1_data = qs_queue_1_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_151 = 6'h1 == deq_id ? deq_bits_1_data : deq_bits_0_data; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_2_data = qs_queue_2_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_152 = 6'h2 == deq_id ? deq_bits_2_data : _GEN_151; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_3_data = qs_queue_3_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_153 = 6'h3 == deq_id ? deq_bits_3_data : _GEN_152; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_4_data = qs_queue_4_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_154 = 6'h4 == deq_id ? deq_bits_4_data : _GEN_153; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_5_data = qs_queue_5_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_155 = 6'h5 == deq_id ? deq_bits_5_data : _GEN_154; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_6_data = qs_queue_6_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_156 = 6'h6 == deq_id ? deq_bits_6_data : _GEN_155; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_7_data = qs_queue_7_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_157 = 6'h7 == deq_id ? deq_bits_7_data : _GEN_156; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_8_data = qs_queue_8_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_158 = 6'h8 == deq_id ? deq_bits_8_data : _GEN_157; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_9_data = qs_queue_9_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_159 = 6'h9 == deq_id ? deq_bits_9_data : _GEN_158; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_10_data = qs_queue_10_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_160 = 6'ha == deq_id ? deq_bits_10_data : _GEN_159; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_11_data = qs_queue_11_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_161 = 6'hb == deq_id ? deq_bits_11_data : _GEN_160; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_12_data = qs_queue_12_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_162 = 6'hc == deq_id ? deq_bits_12_data : _GEN_161; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_13_data = qs_queue_13_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_163 = 6'hd == deq_id ? deq_bits_13_data : _GEN_162; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_14_data = qs_queue_14_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_164 = 6'he == deq_id ? deq_bits_14_data : _GEN_163; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_15_data = qs_queue_15_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_165 = 6'hf == deq_id ? deq_bits_15_data : _GEN_164; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_16_data = qs_queue_16_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_166 = 6'h10 == deq_id ? deq_bits_16_data : _GEN_165; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_17_data = qs_queue_17_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_167 = 6'h11 == deq_id ? deq_bits_17_data : _GEN_166; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_18_data = qs_queue_18_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_168 = 6'h12 == deq_id ? deq_bits_18_data : _GEN_167; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_19_data = qs_queue_19_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_169 = 6'h13 == deq_id ? deq_bits_19_data : _GEN_168; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_20_data = qs_queue_20_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_170 = 6'h14 == deq_id ? deq_bits_20_data : _GEN_169; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_21_data = qs_queue_21_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_171 = 6'h15 == deq_id ? deq_bits_21_data : _GEN_170; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_22_data = qs_queue_22_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_172 = 6'h16 == deq_id ? deq_bits_22_data : _GEN_171; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_23_data = qs_queue_23_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_173 = 6'h17 == deq_id ? deq_bits_23_data : _GEN_172; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_24_data = qs_queue_24_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_174 = 6'h18 == deq_id ? deq_bits_24_data : _GEN_173; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_25_data = qs_queue_25_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_175 = 6'h19 == deq_id ? deq_bits_25_data : _GEN_174; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_26_data = qs_queue_26_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_176 = 6'h1a == deq_id ? deq_bits_26_data : _GEN_175; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_27_data = qs_queue_27_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_177 = 6'h1b == deq_id ? deq_bits_27_data : _GEN_176; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_28_data = qs_queue_28_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_178 = 6'h1c == deq_id ? deq_bits_28_data : _GEN_177; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_29_data = qs_queue_29_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_179 = 6'h1d == deq_id ? deq_bits_29_data : _GEN_178; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_30_data = qs_queue_30_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_180 = 6'h1e == deq_id ? deq_bits_30_data : _GEN_179; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_31_data = qs_queue_31_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_181 = 6'h1f == deq_id ? deq_bits_31_data : _GEN_180; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_32_data = qs_queue_32_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_182 = 6'h20 == deq_id ? deq_bits_32_data : _GEN_181; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_33_data = qs_queue_33_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_183 = 6'h21 == deq_id ? deq_bits_33_data : _GEN_182; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_34_data = qs_queue_34_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_184 = 6'h22 == deq_id ? deq_bits_34_data : _GEN_183; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_35_data = qs_queue_35_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [255:0] _GEN_185 = 6'h23 == deq_id ? deq_bits_35_data : _GEN_184; // @[Deinterleaver.scala 115:{20,20}]
  wire [255:0] deq_bits_36_data = qs_queue_36_io_deq_bits_data; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] deq_bits_0_id = qs_queue_0_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] deq_bits_1_id = qs_queue_1_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_188 = 6'h1 == deq_id ? deq_bits_1_id : deq_bits_0_id; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_2_id = qs_queue_2_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_189 = 6'h2 == deq_id ? deq_bits_2_id : _GEN_188; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_3_id = qs_queue_3_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_190 = 6'h3 == deq_id ? deq_bits_3_id : _GEN_189; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_4_id = qs_queue_4_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_191 = 6'h4 == deq_id ? deq_bits_4_id : _GEN_190; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_5_id = qs_queue_5_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_192 = 6'h5 == deq_id ? deq_bits_5_id : _GEN_191; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_6_id = qs_queue_6_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_193 = 6'h6 == deq_id ? deq_bits_6_id : _GEN_192; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_7_id = qs_queue_7_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_194 = 6'h7 == deq_id ? deq_bits_7_id : _GEN_193; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_8_id = qs_queue_8_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_195 = 6'h8 == deq_id ? deq_bits_8_id : _GEN_194; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_9_id = qs_queue_9_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_196 = 6'h9 == deq_id ? deq_bits_9_id : _GEN_195; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_10_id = qs_queue_10_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_197 = 6'ha == deq_id ? deq_bits_10_id : _GEN_196; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_11_id = qs_queue_11_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_198 = 6'hb == deq_id ? deq_bits_11_id : _GEN_197; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_12_id = qs_queue_12_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_199 = 6'hc == deq_id ? deq_bits_12_id : _GEN_198; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_13_id = qs_queue_13_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_200 = 6'hd == deq_id ? deq_bits_13_id : _GEN_199; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_14_id = qs_queue_14_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_201 = 6'he == deq_id ? deq_bits_14_id : _GEN_200; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_15_id = qs_queue_15_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_202 = 6'hf == deq_id ? deq_bits_15_id : _GEN_201; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_16_id = qs_queue_16_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_203 = 6'h10 == deq_id ? deq_bits_16_id : _GEN_202; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_17_id = qs_queue_17_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_204 = 6'h11 == deq_id ? deq_bits_17_id : _GEN_203; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_18_id = qs_queue_18_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_205 = 6'h12 == deq_id ? deq_bits_18_id : _GEN_204; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_19_id = qs_queue_19_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_206 = 6'h13 == deq_id ? deq_bits_19_id : _GEN_205; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_20_id = qs_queue_20_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_207 = 6'h14 == deq_id ? deq_bits_20_id : _GEN_206; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_21_id = qs_queue_21_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_208 = 6'h15 == deq_id ? deq_bits_21_id : _GEN_207; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_22_id = qs_queue_22_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_209 = 6'h16 == deq_id ? deq_bits_22_id : _GEN_208; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_23_id = qs_queue_23_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_210 = 6'h17 == deq_id ? deq_bits_23_id : _GEN_209; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_24_id = qs_queue_24_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_211 = 6'h18 == deq_id ? deq_bits_24_id : _GEN_210; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_25_id = qs_queue_25_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_212 = 6'h19 == deq_id ? deq_bits_25_id : _GEN_211; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_26_id = qs_queue_26_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_213 = 6'h1a == deq_id ? deq_bits_26_id : _GEN_212; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_27_id = qs_queue_27_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_214 = 6'h1b == deq_id ? deq_bits_27_id : _GEN_213; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_28_id = qs_queue_28_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_215 = 6'h1c == deq_id ? deq_bits_28_id : _GEN_214; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_29_id = qs_queue_29_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_216 = 6'h1d == deq_id ? deq_bits_29_id : _GEN_215; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_30_id = qs_queue_30_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_217 = 6'h1e == deq_id ? deq_bits_30_id : _GEN_216; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_31_id = qs_queue_31_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_218 = 6'h1f == deq_id ? deq_bits_31_id : _GEN_217; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_32_id = qs_queue_32_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_219 = 6'h20 == deq_id ? deq_bits_32_id : _GEN_218; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_33_id = qs_queue_33_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_220 = 6'h21 == deq_id ? deq_bits_33_id : _GEN_219; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_34_id = qs_queue_34_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_221 = 6'h22 == deq_id ? deq_bits_34_id : _GEN_220; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_35_id = qs_queue_35_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  wire [5:0] _GEN_222 = 6'h23 == deq_id ? deq_bits_35_id : _GEN_221; // @[Deinterleaver.scala 115:{20,20}]
  wire [5:0] deq_bits_36_id = qs_queue_36_io_deq_bits_id; // @[Deinterleaver.scala 114:{31,31}]
  Queue_27 qs_queue_0 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_0_clock),
    .reset(qs_queue_0_reset),
    .io_enq_ready(qs_queue_0_io_enq_ready),
    .io_enq_valid(qs_queue_0_io_enq_valid),
    .io_enq_bits_id(qs_queue_0_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_0_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_0_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_0_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_0_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_0_io_enq_bits_last),
    .io_deq_ready(qs_queue_0_io_deq_ready),
    .io_deq_valid(qs_queue_0_io_deq_valid),
    .io_deq_bits_id(qs_queue_0_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_0_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_0_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_0_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_0_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_0_io_deq_bits_last)
  );
  Queue_27 qs_queue_1 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_1_clock),
    .reset(qs_queue_1_reset),
    .io_enq_ready(qs_queue_1_io_enq_ready),
    .io_enq_valid(qs_queue_1_io_enq_valid),
    .io_enq_bits_id(qs_queue_1_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_1_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_1_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_1_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_1_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_1_io_enq_bits_last),
    .io_deq_ready(qs_queue_1_io_deq_ready),
    .io_deq_valid(qs_queue_1_io_deq_valid),
    .io_deq_bits_id(qs_queue_1_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_1_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_1_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_1_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_1_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_1_io_deq_bits_last)
  );
  Queue_27 qs_queue_2 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_2_clock),
    .reset(qs_queue_2_reset),
    .io_enq_ready(qs_queue_2_io_enq_ready),
    .io_enq_valid(qs_queue_2_io_enq_valid),
    .io_enq_bits_id(qs_queue_2_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_2_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_2_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_2_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_2_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_2_io_enq_bits_last),
    .io_deq_ready(qs_queue_2_io_deq_ready),
    .io_deq_valid(qs_queue_2_io_deq_valid),
    .io_deq_bits_id(qs_queue_2_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_2_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_2_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_2_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_2_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_2_io_deq_bits_last)
  );
  Queue_27 qs_queue_3 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_3_clock),
    .reset(qs_queue_3_reset),
    .io_enq_ready(qs_queue_3_io_enq_ready),
    .io_enq_valid(qs_queue_3_io_enq_valid),
    .io_enq_bits_id(qs_queue_3_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_3_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_3_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_3_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_3_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_3_io_enq_bits_last),
    .io_deq_ready(qs_queue_3_io_deq_ready),
    .io_deq_valid(qs_queue_3_io_deq_valid),
    .io_deq_bits_id(qs_queue_3_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_3_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_3_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_3_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_3_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_3_io_deq_bits_last)
  );
  Queue_27 qs_queue_4 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_4_clock),
    .reset(qs_queue_4_reset),
    .io_enq_ready(qs_queue_4_io_enq_ready),
    .io_enq_valid(qs_queue_4_io_enq_valid),
    .io_enq_bits_id(qs_queue_4_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_4_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_4_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_4_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_4_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_4_io_enq_bits_last),
    .io_deq_ready(qs_queue_4_io_deq_ready),
    .io_deq_valid(qs_queue_4_io_deq_valid),
    .io_deq_bits_id(qs_queue_4_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_4_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_4_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_4_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_4_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_4_io_deq_bits_last)
  );
  Queue_27 qs_queue_5 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_5_clock),
    .reset(qs_queue_5_reset),
    .io_enq_ready(qs_queue_5_io_enq_ready),
    .io_enq_valid(qs_queue_5_io_enq_valid),
    .io_enq_bits_id(qs_queue_5_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_5_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_5_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_5_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_5_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_5_io_enq_bits_last),
    .io_deq_ready(qs_queue_5_io_deq_ready),
    .io_deq_valid(qs_queue_5_io_deq_valid),
    .io_deq_bits_id(qs_queue_5_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_5_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_5_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_5_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_5_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_5_io_deq_bits_last)
  );
  Queue_27 qs_queue_6 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_6_clock),
    .reset(qs_queue_6_reset),
    .io_enq_ready(qs_queue_6_io_enq_ready),
    .io_enq_valid(qs_queue_6_io_enq_valid),
    .io_enq_bits_id(qs_queue_6_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_6_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_6_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_6_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_6_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_6_io_enq_bits_last),
    .io_deq_ready(qs_queue_6_io_deq_ready),
    .io_deq_valid(qs_queue_6_io_deq_valid),
    .io_deq_bits_id(qs_queue_6_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_6_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_6_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_6_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_6_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_6_io_deq_bits_last)
  );
  Queue_27 qs_queue_7 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_7_clock),
    .reset(qs_queue_7_reset),
    .io_enq_ready(qs_queue_7_io_enq_ready),
    .io_enq_valid(qs_queue_7_io_enq_valid),
    .io_enq_bits_id(qs_queue_7_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_7_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_7_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_7_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_7_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_7_io_enq_bits_last),
    .io_deq_ready(qs_queue_7_io_deq_ready),
    .io_deq_valid(qs_queue_7_io_deq_valid),
    .io_deq_bits_id(qs_queue_7_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_7_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_7_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_7_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_7_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_7_io_deq_bits_last)
  );
  Queue_27 qs_queue_8 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_8_clock),
    .reset(qs_queue_8_reset),
    .io_enq_ready(qs_queue_8_io_enq_ready),
    .io_enq_valid(qs_queue_8_io_enq_valid),
    .io_enq_bits_id(qs_queue_8_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_8_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_8_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_8_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_8_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_8_io_enq_bits_last),
    .io_deq_ready(qs_queue_8_io_deq_ready),
    .io_deq_valid(qs_queue_8_io_deq_valid),
    .io_deq_bits_id(qs_queue_8_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_8_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_8_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_8_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_8_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_8_io_deq_bits_last)
  );
  Queue_27 qs_queue_9 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_9_clock),
    .reset(qs_queue_9_reset),
    .io_enq_ready(qs_queue_9_io_enq_ready),
    .io_enq_valid(qs_queue_9_io_enq_valid),
    .io_enq_bits_id(qs_queue_9_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_9_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_9_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_9_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_9_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_9_io_enq_bits_last),
    .io_deq_ready(qs_queue_9_io_deq_ready),
    .io_deq_valid(qs_queue_9_io_deq_valid),
    .io_deq_bits_id(qs_queue_9_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_9_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_9_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_9_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_9_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_9_io_deq_bits_last)
  );
  Queue_27 qs_queue_10 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_10_clock),
    .reset(qs_queue_10_reset),
    .io_enq_ready(qs_queue_10_io_enq_ready),
    .io_enq_valid(qs_queue_10_io_enq_valid),
    .io_enq_bits_id(qs_queue_10_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_10_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_10_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_10_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_10_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_10_io_enq_bits_last),
    .io_deq_ready(qs_queue_10_io_deq_ready),
    .io_deq_valid(qs_queue_10_io_deq_valid),
    .io_deq_bits_id(qs_queue_10_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_10_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_10_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_10_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_10_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_10_io_deq_bits_last)
  );
  Queue_27 qs_queue_11 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_11_clock),
    .reset(qs_queue_11_reset),
    .io_enq_ready(qs_queue_11_io_enq_ready),
    .io_enq_valid(qs_queue_11_io_enq_valid),
    .io_enq_bits_id(qs_queue_11_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_11_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_11_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_11_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_11_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_11_io_enq_bits_last),
    .io_deq_ready(qs_queue_11_io_deq_ready),
    .io_deq_valid(qs_queue_11_io_deq_valid),
    .io_deq_bits_id(qs_queue_11_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_11_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_11_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_11_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_11_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_11_io_deq_bits_last)
  );
  Queue_27 qs_queue_12 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_12_clock),
    .reset(qs_queue_12_reset),
    .io_enq_ready(qs_queue_12_io_enq_ready),
    .io_enq_valid(qs_queue_12_io_enq_valid),
    .io_enq_bits_id(qs_queue_12_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_12_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_12_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_12_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_12_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_12_io_enq_bits_last),
    .io_deq_ready(qs_queue_12_io_deq_ready),
    .io_deq_valid(qs_queue_12_io_deq_valid),
    .io_deq_bits_id(qs_queue_12_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_12_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_12_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_12_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_12_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_12_io_deq_bits_last)
  );
  Queue_27 qs_queue_13 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_13_clock),
    .reset(qs_queue_13_reset),
    .io_enq_ready(qs_queue_13_io_enq_ready),
    .io_enq_valid(qs_queue_13_io_enq_valid),
    .io_enq_bits_id(qs_queue_13_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_13_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_13_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_13_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_13_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_13_io_enq_bits_last),
    .io_deq_ready(qs_queue_13_io_deq_ready),
    .io_deq_valid(qs_queue_13_io_deq_valid),
    .io_deq_bits_id(qs_queue_13_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_13_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_13_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_13_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_13_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_13_io_deq_bits_last)
  );
  Queue_27 qs_queue_14 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_14_clock),
    .reset(qs_queue_14_reset),
    .io_enq_ready(qs_queue_14_io_enq_ready),
    .io_enq_valid(qs_queue_14_io_enq_valid),
    .io_enq_bits_id(qs_queue_14_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_14_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_14_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_14_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_14_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_14_io_enq_bits_last),
    .io_deq_ready(qs_queue_14_io_deq_ready),
    .io_deq_valid(qs_queue_14_io_deq_valid),
    .io_deq_bits_id(qs_queue_14_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_14_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_14_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_14_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_14_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_14_io_deq_bits_last)
  );
  Queue_27 qs_queue_15 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_15_clock),
    .reset(qs_queue_15_reset),
    .io_enq_ready(qs_queue_15_io_enq_ready),
    .io_enq_valid(qs_queue_15_io_enq_valid),
    .io_enq_bits_id(qs_queue_15_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_15_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_15_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_15_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_15_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_15_io_enq_bits_last),
    .io_deq_ready(qs_queue_15_io_deq_ready),
    .io_deq_valid(qs_queue_15_io_deq_valid),
    .io_deq_bits_id(qs_queue_15_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_15_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_15_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_15_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_15_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_15_io_deq_bits_last)
  );
  Queue_27 qs_queue_16 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_16_clock),
    .reset(qs_queue_16_reset),
    .io_enq_ready(qs_queue_16_io_enq_ready),
    .io_enq_valid(qs_queue_16_io_enq_valid),
    .io_enq_bits_id(qs_queue_16_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_16_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_16_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_16_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_16_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_16_io_enq_bits_last),
    .io_deq_ready(qs_queue_16_io_deq_ready),
    .io_deq_valid(qs_queue_16_io_deq_valid),
    .io_deq_bits_id(qs_queue_16_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_16_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_16_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_16_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_16_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_16_io_deq_bits_last)
  );
  Queue_27 qs_queue_17 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_17_clock),
    .reset(qs_queue_17_reset),
    .io_enq_ready(qs_queue_17_io_enq_ready),
    .io_enq_valid(qs_queue_17_io_enq_valid),
    .io_enq_bits_id(qs_queue_17_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_17_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_17_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_17_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_17_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_17_io_enq_bits_last),
    .io_deq_ready(qs_queue_17_io_deq_ready),
    .io_deq_valid(qs_queue_17_io_deq_valid),
    .io_deq_bits_id(qs_queue_17_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_17_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_17_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_17_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_17_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_17_io_deq_bits_last)
  );
  Queue_27 qs_queue_18 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_18_clock),
    .reset(qs_queue_18_reset),
    .io_enq_ready(qs_queue_18_io_enq_ready),
    .io_enq_valid(qs_queue_18_io_enq_valid),
    .io_enq_bits_id(qs_queue_18_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_18_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_18_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_18_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_18_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_18_io_enq_bits_last),
    .io_deq_ready(qs_queue_18_io_deq_ready),
    .io_deq_valid(qs_queue_18_io_deq_valid),
    .io_deq_bits_id(qs_queue_18_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_18_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_18_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_18_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_18_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_18_io_deq_bits_last)
  );
  Queue_27 qs_queue_19 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_19_clock),
    .reset(qs_queue_19_reset),
    .io_enq_ready(qs_queue_19_io_enq_ready),
    .io_enq_valid(qs_queue_19_io_enq_valid),
    .io_enq_bits_id(qs_queue_19_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_19_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_19_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_19_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_19_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_19_io_enq_bits_last),
    .io_deq_ready(qs_queue_19_io_deq_ready),
    .io_deq_valid(qs_queue_19_io_deq_valid),
    .io_deq_bits_id(qs_queue_19_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_19_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_19_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_19_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_19_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_19_io_deq_bits_last)
  );
  Queue_27 qs_queue_20 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_20_clock),
    .reset(qs_queue_20_reset),
    .io_enq_ready(qs_queue_20_io_enq_ready),
    .io_enq_valid(qs_queue_20_io_enq_valid),
    .io_enq_bits_id(qs_queue_20_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_20_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_20_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_20_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_20_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_20_io_enq_bits_last),
    .io_deq_ready(qs_queue_20_io_deq_ready),
    .io_deq_valid(qs_queue_20_io_deq_valid),
    .io_deq_bits_id(qs_queue_20_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_20_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_20_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_20_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_20_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_20_io_deq_bits_last)
  );
  Queue_27 qs_queue_21 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_21_clock),
    .reset(qs_queue_21_reset),
    .io_enq_ready(qs_queue_21_io_enq_ready),
    .io_enq_valid(qs_queue_21_io_enq_valid),
    .io_enq_bits_id(qs_queue_21_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_21_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_21_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_21_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_21_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_21_io_enq_bits_last),
    .io_deq_ready(qs_queue_21_io_deq_ready),
    .io_deq_valid(qs_queue_21_io_deq_valid),
    .io_deq_bits_id(qs_queue_21_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_21_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_21_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_21_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_21_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_21_io_deq_bits_last)
  );
  Queue_27 qs_queue_22 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_22_clock),
    .reset(qs_queue_22_reset),
    .io_enq_ready(qs_queue_22_io_enq_ready),
    .io_enq_valid(qs_queue_22_io_enq_valid),
    .io_enq_bits_id(qs_queue_22_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_22_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_22_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_22_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_22_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_22_io_enq_bits_last),
    .io_deq_ready(qs_queue_22_io_deq_ready),
    .io_deq_valid(qs_queue_22_io_deq_valid),
    .io_deq_bits_id(qs_queue_22_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_22_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_22_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_22_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_22_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_22_io_deq_bits_last)
  );
  Queue_27 qs_queue_23 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_23_clock),
    .reset(qs_queue_23_reset),
    .io_enq_ready(qs_queue_23_io_enq_ready),
    .io_enq_valid(qs_queue_23_io_enq_valid),
    .io_enq_bits_id(qs_queue_23_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_23_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_23_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_23_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_23_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_23_io_enq_bits_last),
    .io_deq_ready(qs_queue_23_io_deq_ready),
    .io_deq_valid(qs_queue_23_io_deq_valid),
    .io_deq_bits_id(qs_queue_23_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_23_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_23_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_23_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_23_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_23_io_deq_bits_last)
  );
  Queue_27 qs_queue_24 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_24_clock),
    .reset(qs_queue_24_reset),
    .io_enq_ready(qs_queue_24_io_enq_ready),
    .io_enq_valid(qs_queue_24_io_enq_valid),
    .io_enq_bits_id(qs_queue_24_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_24_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_24_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_24_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_24_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_24_io_enq_bits_last),
    .io_deq_ready(qs_queue_24_io_deq_ready),
    .io_deq_valid(qs_queue_24_io_deq_valid),
    .io_deq_bits_id(qs_queue_24_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_24_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_24_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_24_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_24_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_24_io_deq_bits_last)
  );
  Queue_27 qs_queue_25 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_25_clock),
    .reset(qs_queue_25_reset),
    .io_enq_ready(qs_queue_25_io_enq_ready),
    .io_enq_valid(qs_queue_25_io_enq_valid),
    .io_enq_bits_id(qs_queue_25_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_25_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_25_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_25_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_25_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_25_io_enq_bits_last),
    .io_deq_ready(qs_queue_25_io_deq_ready),
    .io_deq_valid(qs_queue_25_io_deq_valid),
    .io_deq_bits_id(qs_queue_25_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_25_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_25_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_25_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_25_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_25_io_deq_bits_last)
  );
  Queue_27 qs_queue_26 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_26_clock),
    .reset(qs_queue_26_reset),
    .io_enq_ready(qs_queue_26_io_enq_ready),
    .io_enq_valid(qs_queue_26_io_enq_valid),
    .io_enq_bits_id(qs_queue_26_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_26_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_26_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_26_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_26_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_26_io_enq_bits_last),
    .io_deq_ready(qs_queue_26_io_deq_ready),
    .io_deq_valid(qs_queue_26_io_deq_valid),
    .io_deq_bits_id(qs_queue_26_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_26_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_26_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_26_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_26_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_26_io_deq_bits_last)
  );
  Queue_27 qs_queue_27 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_27_clock),
    .reset(qs_queue_27_reset),
    .io_enq_ready(qs_queue_27_io_enq_ready),
    .io_enq_valid(qs_queue_27_io_enq_valid),
    .io_enq_bits_id(qs_queue_27_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_27_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_27_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_27_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_27_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_27_io_enq_bits_last),
    .io_deq_ready(qs_queue_27_io_deq_ready),
    .io_deq_valid(qs_queue_27_io_deq_valid),
    .io_deq_bits_id(qs_queue_27_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_27_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_27_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_27_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_27_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_27_io_deq_bits_last)
  );
  Queue_27 qs_queue_28 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_28_clock),
    .reset(qs_queue_28_reset),
    .io_enq_ready(qs_queue_28_io_enq_ready),
    .io_enq_valid(qs_queue_28_io_enq_valid),
    .io_enq_bits_id(qs_queue_28_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_28_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_28_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_28_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_28_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_28_io_enq_bits_last),
    .io_deq_ready(qs_queue_28_io_deq_ready),
    .io_deq_valid(qs_queue_28_io_deq_valid),
    .io_deq_bits_id(qs_queue_28_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_28_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_28_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_28_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_28_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_28_io_deq_bits_last)
  );
  Queue_27 qs_queue_29 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_29_clock),
    .reset(qs_queue_29_reset),
    .io_enq_ready(qs_queue_29_io_enq_ready),
    .io_enq_valid(qs_queue_29_io_enq_valid),
    .io_enq_bits_id(qs_queue_29_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_29_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_29_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_29_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_29_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_29_io_enq_bits_last),
    .io_deq_ready(qs_queue_29_io_deq_ready),
    .io_deq_valid(qs_queue_29_io_deq_valid),
    .io_deq_bits_id(qs_queue_29_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_29_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_29_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_29_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_29_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_29_io_deq_bits_last)
  );
  Queue_27 qs_queue_30 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_30_clock),
    .reset(qs_queue_30_reset),
    .io_enq_ready(qs_queue_30_io_enq_ready),
    .io_enq_valid(qs_queue_30_io_enq_valid),
    .io_enq_bits_id(qs_queue_30_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_30_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_30_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_30_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_30_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_30_io_enq_bits_last),
    .io_deq_ready(qs_queue_30_io_deq_ready),
    .io_deq_valid(qs_queue_30_io_deq_valid),
    .io_deq_bits_id(qs_queue_30_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_30_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_30_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_30_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_30_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_30_io_deq_bits_last)
  );
  Queue_27 qs_queue_31 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_31_clock),
    .reset(qs_queue_31_reset),
    .io_enq_ready(qs_queue_31_io_enq_ready),
    .io_enq_valid(qs_queue_31_io_enq_valid),
    .io_enq_bits_id(qs_queue_31_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_31_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_31_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_31_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_31_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_31_io_enq_bits_last),
    .io_deq_ready(qs_queue_31_io_deq_ready),
    .io_deq_valid(qs_queue_31_io_deq_valid),
    .io_deq_bits_id(qs_queue_31_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_31_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_31_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_31_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_31_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_31_io_deq_bits_last)
  );
  Queue_27 qs_queue_32 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_32_clock),
    .reset(qs_queue_32_reset),
    .io_enq_ready(qs_queue_32_io_enq_ready),
    .io_enq_valid(qs_queue_32_io_enq_valid),
    .io_enq_bits_id(qs_queue_32_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_32_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_32_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_32_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_32_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_32_io_enq_bits_last),
    .io_deq_ready(qs_queue_32_io_deq_ready),
    .io_deq_valid(qs_queue_32_io_deq_valid),
    .io_deq_bits_id(qs_queue_32_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_32_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_32_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_32_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_32_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_32_io_deq_bits_last)
  );
  Queue_27 qs_queue_33 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_33_clock),
    .reset(qs_queue_33_reset),
    .io_enq_ready(qs_queue_33_io_enq_ready),
    .io_enq_valid(qs_queue_33_io_enq_valid),
    .io_enq_bits_id(qs_queue_33_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_33_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_33_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_33_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_33_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_33_io_enq_bits_last),
    .io_deq_ready(qs_queue_33_io_deq_ready),
    .io_deq_valid(qs_queue_33_io_deq_valid),
    .io_deq_bits_id(qs_queue_33_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_33_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_33_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_33_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_33_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_33_io_deq_bits_last)
  );
  Queue_27 qs_queue_34 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_34_clock),
    .reset(qs_queue_34_reset),
    .io_enq_ready(qs_queue_34_io_enq_ready),
    .io_enq_valid(qs_queue_34_io_enq_valid),
    .io_enq_bits_id(qs_queue_34_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_34_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_34_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_34_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_34_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_34_io_enq_bits_last),
    .io_deq_ready(qs_queue_34_io_deq_ready),
    .io_deq_valid(qs_queue_34_io_deq_valid),
    .io_deq_bits_id(qs_queue_34_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_34_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_34_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_34_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_34_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_34_io_deq_bits_last)
  );
  Queue_27 qs_queue_35 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_35_clock),
    .reset(qs_queue_35_reset),
    .io_enq_ready(qs_queue_35_io_enq_ready),
    .io_enq_valid(qs_queue_35_io_enq_valid),
    .io_enq_bits_id(qs_queue_35_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_35_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_35_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_35_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_35_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_35_io_enq_bits_last),
    .io_deq_ready(qs_queue_35_io_deq_ready),
    .io_deq_valid(qs_queue_35_io_deq_valid),
    .io_deq_bits_id(qs_queue_35_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_35_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_35_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_35_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_35_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_35_io_deq_bits_last)
  );
  Queue_27 qs_queue_36 ( // @[Deinterleaver.scala 66:27]
    .clock(qs_queue_36_clock),
    .reset(qs_queue_36_reset),
    .io_enq_ready(qs_queue_36_io_enq_ready),
    .io_enq_valid(qs_queue_36_io_enq_valid),
    .io_enq_bits_id(qs_queue_36_io_enq_bits_id),
    .io_enq_bits_data(qs_queue_36_io_enq_bits_data),
    .io_enq_bits_resp(qs_queue_36_io_enq_bits_resp),
    .io_enq_bits_echo_tl_state_size(qs_queue_36_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(qs_queue_36_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_last(qs_queue_36_io_enq_bits_last),
    .io_deq_ready(qs_queue_36_io_deq_ready),
    .io_deq_valid(qs_queue_36_io_deq_valid),
    .io_deq_bits_id(qs_queue_36_io_deq_bits_id),
    .io_deq_bits_data(qs_queue_36_io_deq_bits_data),
    .io_deq_bits_resp(qs_queue_36_io_deq_bits_resp),
    .io_deq_bits_echo_tl_state_size(qs_queue_36_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(qs_queue_36_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_last(qs_queue_36_io_deq_bits_last)
  );
  assign auto_in_awready = auto_out_awready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_wready = auto_out_wready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bvalid = auto_out_bvalid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bid = auto_out_bid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_bresp = auto_out_bresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_becho_tl_state_size = auto_out_becho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_becho_tl_state_source = auto_out_becho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_arready = auto_out_arready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign auto_in_rvalid = locked; // @[Deinterleaver.scala 113:20 Nodes.scala 1210:84]
  assign auto_in_rid = 6'h24 == deq_id ? deq_bits_36_id : _GEN_222; // @[Deinterleaver.scala 115:{20,20}]
  assign auto_in_rdata = 6'h24 == deq_id ? deq_bits_36_data : _GEN_185; // @[Deinterleaver.scala 115:{20,20}]
  assign auto_in_rresp = 6'h24 == deq_id ? deq_bits_36_resp : _GEN_148; // @[Deinterleaver.scala 115:{20,20}]
  assign auto_in_recho_tl_state_size = 6'h24 == deq_id ? deq_bits_36_echo_tl_state_size : _GEN_111; // @[Deinterleaver.scala 115:{20,20}]
  assign auto_in_recho_tl_state_source = 6'h24 == deq_id ? deq_bits_36_echo_tl_state_source : _GEN_74; // @[Deinterleaver.scala 115:{20,20}]
  assign auto_in_rlast = 6'h24 == deq_id ? deq_bits_36_last : _GEN_37; // @[Deinterleaver.scala 115:{20,20}]
  assign auto_out_awvalid = auto_in_awvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awid = auto_in_awid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awaddr = auto_in_awaddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awlen = auto_in_awlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awsize = auto_in_awsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awburst = auto_in_awburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awlock = auto_in_awlock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awcache = auto_in_awcache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awprot = auto_in_awprot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awqos = auto_in_awqos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awecho_tl_state_size = auto_in_awecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_awecho_tl_state_source = auto_in_awecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wvalid = auto_in_wvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wdata = auto_in_wdata; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wstrb = auto_in_wstrb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_wlast = auto_in_wlast; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_bready = auto_in_bready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arvalid = auto_in_arvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arid = auto_in_arid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_araddr = auto_in_araddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arlen = auto_in_arlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arsize = auto_in_arsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arburst = auto_in_arburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arlock = auto_in_arlock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arcache = auto_in_arcache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arprot = auto_in_arprot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arqos = auto_in_arqos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arecho_tl_state_size = auto_in_arecho_tl_state_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_arecho_tl_state_source = auto_in_arecho_tl_state_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign auto_out_rready = 6'h24 == auto_out_rid ? enq_readys_36 : _GEN_259; // @[Deinterleaver.scala 126:{21,21}]
  assign qs_queue_0_clock = clock;
  assign qs_queue_0_reset = reset;
  assign qs_queue_0_io_enq_valid = enq_OH[0] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_0_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_0_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_0_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_0_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_0_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_0_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_0_io_deq_ready = deq_OH[0] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_1_clock = clock;
  assign qs_queue_1_reset = reset;
  assign qs_queue_1_io_enq_valid = enq_OH[1] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_1_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_1_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_1_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_1_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_1_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_1_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_1_io_deq_ready = deq_OH[1] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_2_clock = clock;
  assign qs_queue_2_reset = reset;
  assign qs_queue_2_io_enq_valid = enq_OH[2] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_2_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_2_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_2_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_2_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_2_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_2_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_2_io_deq_ready = deq_OH[2] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_3_clock = clock;
  assign qs_queue_3_reset = reset;
  assign qs_queue_3_io_enq_valid = enq_OH[3] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_3_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_3_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_3_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_3_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_3_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_3_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_3_io_deq_ready = deq_OH[3] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_4_clock = clock;
  assign qs_queue_4_reset = reset;
  assign qs_queue_4_io_enq_valid = enq_OH[4] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_4_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_4_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_4_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_4_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_4_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_4_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_4_io_deq_ready = deq_OH[4] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_5_clock = clock;
  assign qs_queue_5_reset = reset;
  assign qs_queue_5_io_enq_valid = enq_OH[5] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_5_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_5_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_5_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_5_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_5_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_5_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_5_io_deq_ready = deq_OH[5] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_6_clock = clock;
  assign qs_queue_6_reset = reset;
  assign qs_queue_6_io_enq_valid = enq_OH[6] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_6_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_6_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_6_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_6_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_6_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_6_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_6_io_deq_ready = deq_OH[6] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_7_clock = clock;
  assign qs_queue_7_reset = reset;
  assign qs_queue_7_io_enq_valid = enq_OH[7] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_7_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_7_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_7_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_7_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_7_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_7_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_7_io_deq_ready = deq_OH[7] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_8_clock = clock;
  assign qs_queue_8_reset = reset;
  assign qs_queue_8_io_enq_valid = enq_OH[8] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_8_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_8_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_8_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_8_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_8_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_8_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_8_io_deq_ready = deq_OH[8] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_9_clock = clock;
  assign qs_queue_9_reset = reset;
  assign qs_queue_9_io_enq_valid = enq_OH[9] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_9_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_9_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_9_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_9_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_9_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_9_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_9_io_deq_ready = deq_OH[9] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_10_clock = clock;
  assign qs_queue_10_reset = reset;
  assign qs_queue_10_io_enq_valid = enq_OH[10] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_10_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_10_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_10_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_10_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_10_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_10_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_10_io_deq_ready = deq_OH[10] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_11_clock = clock;
  assign qs_queue_11_reset = reset;
  assign qs_queue_11_io_enq_valid = enq_OH[11] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_11_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_11_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_11_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_11_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_11_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_11_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_11_io_deq_ready = deq_OH[11] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_12_clock = clock;
  assign qs_queue_12_reset = reset;
  assign qs_queue_12_io_enq_valid = enq_OH[12] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_12_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_12_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_12_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_12_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_12_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_12_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_12_io_deq_ready = deq_OH[12] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_13_clock = clock;
  assign qs_queue_13_reset = reset;
  assign qs_queue_13_io_enq_valid = enq_OH[13] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_13_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_13_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_13_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_13_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_13_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_13_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_13_io_deq_ready = deq_OH[13] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_14_clock = clock;
  assign qs_queue_14_reset = reset;
  assign qs_queue_14_io_enq_valid = enq_OH[14] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_14_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_14_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_14_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_14_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_14_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_14_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_14_io_deq_ready = deq_OH[14] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_15_clock = clock;
  assign qs_queue_15_reset = reset;
  assign qs_queue_15_io_enq_valid = enq_OH[15] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_15_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_15_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_15_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_15_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_15_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_15_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_15_io_deq_ready = deq_OH[15] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_16_clock = clock;
  assign qs_queue_16_reset = reset;
  assign qs_queue_16_io_enq_valid = enq_OH[16] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_16_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_16_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_16_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_16_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_16_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_16_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_16_io_deq_ready = deq_OH[16] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_17_clock = clock;
  assign qs_queue_17_reset = reset;
  assign qs_queue_17_io_enq_valid = enq_OH[17] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_17_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_17_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_17_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_17_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_17_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_17_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_17_io_deq_ready = deq_OH[17] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_18_clock = clock;
  assign qs_queue_18_reset = reset;
  assign qs_queue_18_io_enq_valid = enq_OH[18] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_18_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_18_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_18_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_18_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_18_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_18_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_18_io_deq_ready = deq_OH[18] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_19_clock = clock;
  assign qs_queue_19_reset = reset;
  assign qs_queue_19_io_enq_valid = enq_OH[19] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_19_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_19_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_19_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_19_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_19_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_19_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_19_io_deq_ready = deq_OH[19] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_20_clock = clock;
  assign qs_queue_20_reset = reset;
  assign qs_queue_20_io_enq_valid = enq_OH[20] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_20_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_20_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_20_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_20_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_20_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_20_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_20_io_deq_ready = deq_OH[20] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_21_clock = clock;
  assign qs_queue_21_reset = reset;
  assign qs_queue_21_io_enq_valid = enq_OH[21] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_21_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_21_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_21_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_21_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_21_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_21_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_21_io_deq_ready = deq_OH[21] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_22_clock = clock;
  assign qs_queue_22_reset = reset;
  assign qs_queue_22_io_enq_valid = enq_OH[22] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_22_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_22_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_22_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_22_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_22_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_22_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_22_io_deq_ready = deq_OH[22] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_23_clock = clock;
  assign qs_queue_23_reset = reset;
  assign qs_queue_23_io_enq_valid = enq_OH[23] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_23_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_23_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_23_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_23_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_23_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_23_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_23_io_deq_ready = deq_OH[23] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_24_clock = clock;
  assign qs_queue_24_reset = reset;
  assign qs_queue_24_io_enq_valid = enq_OH[24] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_24_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_24_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_24_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_24_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_24_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_24_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_24_io_deq_ready = deq_OH[24] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_25_clock = clock;
  assign qs_queue_25_reset = reset;
  assign qs_queue_25_io_enq_valid = enq_OH[25] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_25_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_25_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_25_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_25_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_25_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_25_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_25_io_deq_ready = deq_OH[25] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_26_clock = clock;
  assign qs_queue_26_reset = reset;
  assign qs_queue_26_io_enq_valid = enq_OH[26] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_26_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_26_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_26_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_26_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_26_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_26_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_26_io_deq_ready = deq_OH[26] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_27_clock = clock;
  assign qs_queue_27_reset = reset;
  assign qs_queue_27_io_enq_valid = enq_OH[27] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_27_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_27_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_27_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_27_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_27_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_27_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_27_io_deq_ready = deq_OH[27] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_28_clock = clock;
  assign qs_queue_28_reset = reset;
  assign qs_queue_28_io_enq_valid = enq_OH[28] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_28_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_28_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_28_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_28_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_28_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_28_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_28_io_deq_ready = deq_OH[28] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_29_clock = clock;
  assign qs_queue_29_reset = reset;
  assign qs_queue_29_io_enq_valid = enq_OH[29] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_29_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_29_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_29_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_29_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_29_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_29_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_29_io_deq_ready = deq_OH[29] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_30_clock = clock;
  assign qs_queue_30_reset = reset;
  assign qs_queue_30_io_enq_valid = enq_OH[30] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_30_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_30_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_30_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_30_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_30_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_30_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_30_io_deq_ready = deq_OH[30] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_31_clock = clock;
  assign qs_queue_31_reset = reset;
  assign qs_queue_31_io_enq_valid = enq_OH[31] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_31_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_31_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_31_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_31_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_31_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_31_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_31_io_deq_ready = deq_OH[31] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_32_clock = clock;
  assign qs_queue_32_reset = reset;
  assign qs_queue_32_io_enq_valid = enq_OH[32] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_32_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_32_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_32_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_32_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_32_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_32_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_32_io_deq_ready = deq_OH[32] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_33_clock = clock;
  assign qs_queue_33_reset = reset;
  assign qs_queue_33_io_enq_valid = enq_OH[33] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_33_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_33_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_33_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_33_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_33_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_33_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_33_io_deq_ready = deq_OH[33] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_34_clock = clock;
  assign qs_queue_34_reset = reset;
  assign qs_queue_34_io_enq_valid = enq_OH[34] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_34_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_34_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_34_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_34_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_34_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_34_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_34_io_deq_ready = deq_OH[34] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_35_clock = clock;
  assign qs_queue_35_reset = reset;
  assign qs_queue_35_io_enq_valid = enq_OH[35] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_35_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_35_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_35_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_35_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_35_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_35_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_35_io_deq_ready = deq_OH[35] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  assign qs_queue_36_clock = clock;
  assign qs_queue_36_reset = reset;
  assign qs_queue_36_io_enq_valid = enq_OH[36] & auto_out_rvalid; // @[Deinterleaver.scala 128:28]
  assign qs_queue_36_io_enq_bits_id = auto_out_rid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_36_io_enq_bits_data = auto_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_36_io_enq_bits_resp = auto_out_rresp; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_36_io_enq_bits_echo_tl_state_size = auto_out_recho_tl_state_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_36_io_enq_bits_echo_tl_state_source = auto_out_recho_tl_state_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_36_io_enq_bits_last = auto_out_rlast; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign qs_queue_36_io_deq_ready = deq_OH[36] & _pending_dec_T_1; // @[Deinterleaver.scala 119:28]
  always @(posedge clock) begin
    if (~locked | _pending_dec_T_1 & bundleIn_0_rlast) begin // @[Deinterleaver.scala 107:59]
      deq_id <= _deq_id_T_15; // @[Deinterleaver.scala 109:18]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 107:59]
      locked <= 1'h0; // @[Deinterleaver.scala 108:18]
    end else if (~locked | _pending_dec_T_1 & bundleIn_0_rlast) begin // @[Deinterleaver.scala 82:29]
      locked <= |pending;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count <= 2'h0;
    end else begin
      pending_count <= _pending_next_T_1 - _GEN_262;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_1 <= 2'h0;
    end else begin
      pending_count_1 <= _pending_next_T_5 - _GEN_264;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_2 <= 2'h0;
    end else begin
      pending_count_2 <= _pending_next_T_9 - _GEN_266;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_3 <= 2'h0;
    end else begin
      pending_count_3 <= _pending_next_T_13 - _GEN_268;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_4 <= 2'h0;
    end else begin
      pending_count_4 <= _pending_next_T_17 - _GEN_270;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_5 <= 2'h0;
    end else begin
      pending_count_5 <= _pending_next_T_21 - _GEN_272;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_6 <= 2'h0;
    end else begin
      pending_count_6 <= _pending_next_T_25 - _GEN_274;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_7 <= 2'h0;
    end else begin
      pending_count_7 <= _pending_next_T_29 - _GEN_276;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_8 <= 2'h0;
    end else begin
      pending_count_8 <= _pending_next_T_33 - _GEN_278;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_9 <= 2'h0;
    end else begin
      pending_count_9 <= _pending_next_T_37 - _GEN_280;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_10 <= 2'h0;
    end else begin
      pending_count_10 <= _pending_next_T_41 - _GEN_282;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_11 <= 2'h0;
    end else begin
      pending_count_11 <= _pending_next_T_45 - _GEN_284;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_12 <= 2'h0;
    end else begin
      pending_count_12 <= _pending_next_T_49 - _GEN_286;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_13 <= 2'h0;
    end else begin
      pending_count_13 <= _pending_next_T_53 - _GEN_288;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_14 <= 2'h0;
    end else begin
      pending_count_14 <= _pending_next_T_57 - _GEN_290;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_15 <= 2'h0;
    end else begin
      pending_count_15 <= _pending_next_T_61 - _GEN_292;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_16 <= 2'h0;
    end else begin
      pending_count_16 <= _pending_next_T_65 - _GEN_294;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_17 <= 2'h0;
    end else begin
      pending_count_17 <= _pending_next_T_69 - _GEN_296;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_18 <= 2'h0;
    end else begin
      pending_count_18 <= _pending_next_T_73 - _GEN_298;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_19 <= 2'h0;
    end else begin
      pending_count_19 <= _pending_next_T_77 - _GEN_300;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_20 <= 2'h0;
    end else begin
      pending_count_20 <= _pending_next_T_81 - _GEN_302;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_21 <= 2'h0;
    end else begin
      pending_count_21 <= _pending_next_T_85 - _GEN_304;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_22 <= 2'h0;
    end else begin
      pending_count_22 <= _pending_next_T_89 - _GEN_306;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_23 <= 2'h0;
    end else begin
      pending_count_23 <= _pending_next_T_93 - _GEN_308;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_24 <= 2'h0;
    end else begin
      pending_count_24 <= _pending_next_T_97 - _GEN_310;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_25 <= 2'h0;
    end else begin
      pending_count_25 <= _pending_next_T_101 - _GEN_312;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_26 <= 2'h0;
    end else begin
      pending_count_26 <= _pending_next_T_105 - _GEN_314;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_27 <= 2'h0;
    end else begin
      pending_count_27 <= _pending_next_T_109 - _GEN_316;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_28 <= 2'h0;
    end else begin
      pending_count_28 <= _pending_next_T_113 - _GEN_318;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_29 <= 2'h0;
    end else begin
      pending_count_29 <= _pending_next_T_117 - _GEN_320;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_30 <= 2'h0;
    end else begin
      pending_count_30 <= _pending_next_T_121 - _GEN_322;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_31 <= 2'h0;
    end else begin
      pending_count_31 <= _pending_next_T_125 - _GEN_324;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_32 <= 2'h0;
    end else begin
      pending_count_32 <= _pending_next_T_129 - _GEN_326;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_33 <= 2'h0;
    end else begin
      pending_count_33 <= _pending_next_T_133 - _GEN_328;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_34 <= 2'h0;
    end else begin
      pending_count_34 <= _pending_next_T_137 - _GEN_330;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_35 <= 2'h0;
    end else begin
      pending_count_35 <= _pending_next_T_141 - _GEN_332;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Deinterleaver.scala 96:40]
      pending_count_36 <= 2'h0;
    end else begin
      pending_count_36 <= _pending_next_T_145 - _GEN_334;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  locked = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  deq_id = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  pending_count = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pending_count_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  pending_count_2 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  pending_count_3 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  pending_count_4 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  pending_count_5 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  pending_count_6 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  pending_count_7 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  pending_count_8 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  pending_count_9 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  pending_count_10 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  pending_count_11 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  pending_count_12 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  pending_count_13 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  pending_count_14 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  pending_count_15 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  pending_count_16 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  pending_count_17 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  pending_count_18 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  pending_count_19 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  pending_count_20 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  pending_count_21 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  pending_count_22 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  pending_count_23 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  pending_count_24 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  pending_count_25 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  pending_count_26 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  pending_count_27 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  pending_count_28 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  pending_count_29 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  pending_count_30 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  pending_count_31 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  pending_count_32 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  pending_count_33 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  pending_count_34 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  pending_count_35 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  pending_count_36 = _RAND_38[1:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    locked = 1'h0;
  end
  if (reset) begin
    pending_count = 2'h0;
  end
  if (reset) begin
    pending_count_1 = 2'h0;
  end
  if (reset) begin
    pending_count_2 = 2'h0;
  end
  if (reset) begin
    pending_count_3 = 2'h0;
  end
  if (reset) begin
    pending_count_4 = 2'h0;
  end
  if (reset) begin
    pending_count_5 = 2'h0;
  end
  if (reset) begin
    pending_count_6 = 2'h0;
  end
  if (reset) begin
    pending_count_7 = 2'h0;
  end
  if (reset) begin
    pending_count_8 = 2'h0;
  end
  if (reset) begin
    pending_count_9 = 2'h0;
  end
  if (reset) begin
    pending_count_10 = 2'h0;
  end
  if (reset) begin
    pending_count_11 = 2'h0;
  end
  if (reset) begin
    pending_count_12 = 2'h0;
  end
  if (reset) begin
    pending_count_13 = 2'h0;
  end
  if (reset) begin
    pending_count_14 = 2'h0;
  end
  if (reset) begin
    pending_count_15 = 2'h0;
  end
  if (reset) begin
    pending_count_16 = 2'h0;
  end
  if (reset) begin
    pending_count_17 = 2'h0;
  end
  if (reset) begin
    pending_count_18 = 2'h0;
  end
  if (reset) begin
    pending_count_19 = 2'h0;
  end
  if (reset) begin
    pending_count_20 = 2'h0;
  end
  if (reset) begin
    pending_count_21 = 2'h0;
  end
  if (reset) begin
    pending_count_22 = 2'h0;
  end
  if (reset) begin
    pending_count_23 = 2'h0;
  end
  if (reset) begin
    pending_count_24 = 2'h0;
  end
  if (reset) begin
    pending_count_25 = 2'h0;
  end
  if (reset) begin
    pending_count_26 = 2'h0;
  end
  if (reset) begin
    pending_count_27 = 2'h0;
  end
  if (reset) begin
    pending_count_28 = 2'h0;
  end
  if (reset) begin
    pending_count_29 = 2'h0;
  end
  if (reset) begin
    pending_count_30 = 2'h0;
  end
  if (reset) begin
    pending_count_31 = 2'h0;
  end
  if (reset) begin
    pending_count_32 = 2'h0;
  end
  if (reset) begin
    pending_count_33 = 2'h0;
  end
  if (reset) begin
    pending_count_34 = 2'h0;
  end
  if (reset) begin
    pending_count_35 = 2'h0;
  end
  if (reset) begin
    pending_count_36 = 2'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

