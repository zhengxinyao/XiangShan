module LZA_2(
  input  [48:0] io_a,
  input  [48:0] io_b,
  output [48:0] io_f
);
  wire  k_0 = ~io_a[0] & ~io_b[0]; // @[LZA.scala 19:21]
  wire  p_1 = io_a[1] ^ io_b[1]; // @[LZA.scala 18:18]
  wire  k_1 = ~io_a[1] & ~io_b[1]; // @[LZA.scala 19:21]
  wire  f_1 = p_1 ^ ~k_0; // @[LZA.scala 23:20]
  wire  p_2 = io_a[2] ^ io_b[2]; // @[LZA.scala 18:18]
  wire  k_2 = ~io_a[2] & ~io_b[2]; // @[LZA.scala 19:21]
  wire  f_2 = p_2 ^ ~k_1; // @[LZA.scala 23:20]
  wire  p_3 = io_a[3] ^ io_b[3]; // @[LZA.scala 18:18]
  wire  k_3 = ~io_a[3] & ~io_b[3]; // @[LZA.scala 19:21]
  wire  f_3 = p_3 ^ ~k_2; // @[LZA.scala 23:20]
  wire  p_4 = io_a[4] ^ io_b[4]; // @[LZA.scala 18:18]
  wire  k_4 = ~io_a[4] & ~io_b[4]; // @[LZA.scala 19:21]
  wire  f_4 = p_4 ^ ~k_3; // @[LZA.scala 23:20]
  wire  p_5 = io_a[5] ^ io_b[5]; // @[LZA.scala 18:18]
  wire  k_5 = ~io_a[5] & ~io_b[5]; // @[LZA.scala 19:21]
  wire  f_5 = p_5 ^ ~k_4; // @[LZA.scala 23:20]
  wire  p_6 = io_a[6] ^ io_b[6]; // @[LZA.scala 18:18]
  wire  k_6 = ~io_a[6] & ~io_b[6]; // @[LZA.scala 19:21]
  wire  f_6 = p_6 ^ ~k_5; // @[LZA.scala 23:20]
  wire  p_7 = io_a[7] ^ io_b[7]; // @[LZA.scala 18:18]
  wire  k_7 = ~io_a[7] & ~io_b[7]; // @[LZA.scala 19:21]
  wire  f_7 = p_7 ^ ~k_6; // @[LZA.scala 23:20]
  wire  p_8 = io_a[8] ^ io_b[8]; // @[LZA.scala 18:18]
  wire  k_8 = ~io_a[8] & ~io_b[8]; // @[LZA.scala 19:21]
  wire  f_8 = p_8 ^ ~k_7; // @[LZA.scala 23:20]
  wire  p_9 = io_a[9] ^ io_b[9]; // @[LZA.scala 18:18]
  wire  k_9 = ~io_a[9] & ~io_b[9]; // @[LZA.scala 19:21]
  wire  f_9 = p_9 ^ ~k_8; // @[LZA.scala 23:20]
  wire  p_10 = io_a[10] ^ io_b[10]; // @[LZA.scala 18:18]
  wire  k_10 = ~io_a[10] & ~io_b[10]; // @[LZA.scala 19:21]
  wire  f_10 = p_10 ^ ~k_9; // @[LZA.scala 23:20]
  wire  p_11 = io_a[11] ^ io_b[11]; // @[LZA.scala 18:18]
  wire  k_11 = ~io_a[11] & ~io_b[11]; // @[LZA.scala 19:21]
  wire  f_11 = p_11 ^ ~k_10; // @[LZA.scala 23:20]
  wire  p_12 = io_a[12] ^ io_b[12]; // @[LZA.scala 18:18]
  wire  k_12 = ~io_a[12] & ~io_b[12]; // @[LZA.scala 19:21]
  wire  f_12 = p_12 ^ ~k_11; // @[LZA.scala 23:20]
  wire  p_13 = io_a[13] ^ io_b[13]; // @[LZA.scala 18:18]
  wire  k_13 = ~io_a[13] & ~io_b[13]; // @[LZA.scala 19:21]
  wire  f_13 = p_13 ^ ~k_12; // @[LZA.scala 23:20]
  wire  p_14 = io_a[14] ^ io_b[14]; // @[LZA.scala 18:18]
  wire  k_14 = ~io_a[14] & ~io_b[14]; // @[LZA.scala 19:21]
  wire  f_14 = p_14 ^ ~k_13; // @[LZA.scala 23:20]
  wire  p_15 = io_a[15] ^ io_b[15]; // @[LZA.scala 18:18]
  wire  k_15 = ~io_a[15] & ~io_b[15]; // @[LZA.scala 19:21]
  wire  f_15 = p_15 ^ ~k_14; // @[LZA.scala 23:20]
  wire  p_16 = io_a[16] ^ io_b[16]; // @[LZA.scala 18:18]
  wire  k_16 = ~io_a[16] & ~io_b[16]; // @[LZA.scala 19:21]
  wire  f_16 = p_16 ^ ~k_15; // @[LZA.scala 23:20]
  wire  p_17 = io_a[17] ^ io_b[17]; // @[LZA.scala 18:18]
  wire  k_17 = ~io_a[17] & ~io_b[17]; // @[LZA.scala 19:21]
  wire  f_17 = p_17 ^ ~k_16; // @[LZA.scala 23:20]
  wire  p_18 = io_a[18] ^ io_b[18]; // @[LZA.scala 18:18]
  wire  k_18 = ~io_a[18] & ~io_b[18]; // @[LZA.scala 19:21]
  wire  f_18 = p_18 ^ ~k_17; // @[LZA.scala 23:20]
  wire  p_19 = io_a[19] ^ io_b[19]; // @[LZA.scala 18:18]
  wire  k_19 = ~io_a[19] & ~io_b[19]; // @[LZA.scala 19:21]
  wire  f_19 = p_19 ^ ~k_18; // @[LZA.scala 23:20]
  wire  p_20 = io_a[20] ^ io_b[20]; // @[LZA.scala 18:18]
  wire  k_20 = ~io_a[20] & ~io_b[20]; // @[LZA.scala 19:21]
  wire  f_20 = p_20 ^ ~k_19; // @[LZA.scala 23:20]
  wire  p_21 = io_a[21] ^ io_b[21]; // @[LZA.scala 18:18]
  wire  k_21 = ~io_a[21] & ~io_b[21]; // @[LZA.scala 19:21]
  wire  f_21 = p_21 ^ ~k_20; // @[LZA.scala 23:20]
  wire  p_22 = io_a[22] ^ io_b[22]; // @[LZA.scala 18:18]
  wire  k_22 = ~io_a[22] & ~io_b[22]; // @[LZA.scala 19:21]
  wire  f_22 = p_22 ^ ~k_21; // @[LZA.scala 23:20]
  wire  p_23 = io_a[23] ^ io_b[23]; // @[LZA.scala 18:18]
  wire  k_23 = ~io_a[23] & ~io_b[23]; // @[LZA.scala 19:21]
  wire  f_23 = p_23 ^ ~k_22; // @[LZA.scala 23:20]
  wire  p_24 = io_a[24] ^ io_b[24]; // @[LZA.scala 18:18]
  wire  k_24 = ~io_a[24] & ~io_b[24]; // @[LZA.scala 19:21]
  wire  f_24 = p_24 ^ ~k_23; // @[LZA.scala 23:20]
  wire  p_25 = io_a[25] ^ io_b[25]; // @[LZA.scala 18:18]
  wire  k_25 = ~io_a[25] & ~io_b[25]; // @[LZA.scala 19:21]
  wire  f_25 = p_25 ^ ~k_24; // @[LZA.scala 23:20]
  wire  p_26 = io_a[26] ^ io_b[26]; // @[LZA.scala 18:18]
  wire  k_26 = ~io_a[26] & ~io_b[26]; // @[LZA.scala 19:21]
  wire  f_26 = p_26 ^ ~k_25; // @[LZA.scala 23:20]
  wire  p_27 = io_a[27] ^ io_b[27]; // @[LZA.scala 18:18]
  wire  k_27 = ~io_a[27] & ~io_b[27]; // @[LZA.scala 19:21]
  wire  f_27 = p_27 ^ ~k_26; // @[LZA.scala 23:20]
  wire  p_28 = io_a[28] ^ io_b[28]; // @[LZA.scala 18:18]
  wire  k_28 = ~io_a[28] & ~io_b[28]; // @[LZA.scala 19:21]
  wire  f_28 = p_28 ^ ~k_27; // @[LZA.scala 23:20]
  wire  p_29 = io_a[29] ^ io_b[29]; // @[LZA.scala 18:18]
  wire  k_29 = ~io_a[29] & ~io_b[29]; // @[LZA.scala 19:21]
  wire  f_29 = p_29 ^ ~k_28; // @[LZA.scala 23:20]
  wire  p_30 = io_a[30] ^ io_b[30]; // @[LZA.scala 18:18]
  wire  k_30 = ~io_a[30] & ~io_b[30]; // @[LZA.scala 19:21]
  wire  f_30 = p_30 ^ ~k_29; // @[LZA.scala 23:20]
  wire  p_31 = io_a[31] ^ io_b[31]; // @[LZA.scala 18:18]
  wire  k_31 = ~io_a[31] & ~io_b[31]; // @[LZA.scala 19:21]
  wire  f_31 = p_31 ^ ~k_30; // @[LZA.scala 23:20]
  wire  p_32 = io_a[32] ^ io_b[32]; // @[LZA.scala 18:18]
  wire  k_32 = ~io_a[32] & ~io_b[32]; // @[LZA.scala 19:21]
  wire  f_32 = p_32 ^ ~k_31; // @[LZA.scala 23:20]
  wire  p_33 = io_a[33] ^ io_b[33]; // @[LZA.scala 18:18]
  wire  k_33 = ~io_a[33] & ~io_b[33]; // @[LZA.scala 19:21]
  wire  f_33 = p_33 ^ ~k_32; // @[LZA.scala 23:20]
  wire  p_34 = io_a[34] ^ io_b[34]; // @[LZA.scala 18:18]
  wire  k_34 = ~io_a[34] & ~io_b[34]; // @[LZA.scala 19:21]
  wire  f_34 = p_34 ^ ~k_33; // @[LZA.scala 23:20]
  wire  p_35 = io_a[35] ^ io_b[35]; // @[LZA.scala 18:18]
  wire  k_35 = ~io_a[35] & ~io_b[35]; // @[LZA.scala 19:21]
  wire  f_35 = p_35 ^ ~k_34; // @[LZA.scala 23:20]
  wire  p_36 = io_a[36] ^ io_b[36]; // @[LZA.scala 18:18]
  wire  k_36 = ~io_a[36] & ~io_b[36]; // @[LZA.scala 19:21]
  wire  f_36 = p_36 ^ ~k_35; // @[LZA.scala 23:20]
  wire  p_37 = io_a[37] ^ io_b[37]; // @[LZA.scala 18:18]
  wire  k_37 = ~io_a[37] & ~io_b[37]; // @[LZA.scala 19:21]
  wire  f_37 = p_37 ^ ~k_36; // @[LZA.scala 23:20]
  wire  p_38 = io_a[38] ^ io_b[38]; // @[LZA.scala 18:18]
  wire  k_38 = ~io_a[38] & ~io_b[38]; // @[LZA.scala 19:21]
  wire  f_38 = p_38 ^ ~k_37; // @[LZA.scala 23:20]
  wire  p_39 = io_a[39] ^ io_b[39]; // @[LZA.scala 18:18]
  wire  k_39 = ~io_a[39] & ~io_b[39]; // @[LZA.scala 19:21]
  wire  f_39 = p_39 ^ ~k_38; // @[LZA.scala 23:20]
  wire  p_40 = io_a[40] ^ io_b[40]; // @[LZA.scala 18:18]
  wire  k_40 = ~io_a[40] & ~io_b[40]; // @[LZA.scala 19:21]
  wire  f_40 = p_40 ^ ~k_39; // @[LZA.scala 23:20]
  wire  p_41 = io_a[41] ^ io_b[41]; // @[LZA.scala 18:18]
  wire  k_41 = ~io_a[41] & ~io_b[41]; // @[LZA.scala 19:21]
  wire  f_41 = p_41 ^ ~k_40; // @[LZA.scala 23:20]
  wire  p_42 = io_a[42] ^ io_b[42]; // @[LZA.scala 18:18]
  wire  k_42 = ~io_a[42] & ~io_b[42]; // @[LZA.scala 19:21]
  wire  f_42 = p_42 ^ ~k_41; // @[LZA.scala 23:20]
  wire  p_43 = io_a[43] ^ io_b[43]; // @[LZA.scala 18:18]
  wire  k_43 = ~io_a[43] & ~io_b[43]; // @[LZA.scala 19:21]
  wire  f_43 = p_43 ^ ~k_42; // @[LZA.scala 23:20]
  wire  p_44 = io_a[44] ^ io_b[44]; // @[LZA.scala 18:18]
  wire  k_44 = ~io_a[44] & ~io_b[44]; // @[LZA.scala 19:21]
  wire  f_44 = p_44 ^ ~k_43; // @[LZA.scala 23:20]
  wire  p_45 = io_a[45] ^ io_b[45]; // @[LZA.scala 18:18]
  wire  k_45 = ~io_a[45] & ~io_b[45]; // @[LZA.scala 19:21]
  wire  f_45 = p_45 ^ ~k_44; // @[LZA.scala 23:20]
  wire  p_46 = io_a[46] ^ io_b[46]; // @[LZA.scala 18:18]
  wire  k_46 = ~io_a[46] & ~io_b[46]; // @[LZA.scala 19:21]
  wire  f_46 = p_46 ^ ~k_45; // @[LZA.scala 23:20]
  wire  p_47 = io_a[47] ^ io_b[47]; // @[LZA.scala 18:18]
  wire  k_47 = ~io_a[47] & ~io_b[47]; // @[LZA.scala 19:21]
  wire  f_47 = p_47 ^ ~k_46; // @[LZA.scala 23:20]
  wire  p_48 = io_a[48] ^ io_b[48]; // @[LZA.scala 18:18]
  wire  f_48 = p_48 ^ ~k_47; // @[LZA.scala 23:20]
  wire [5:0] io_f_lo_lo_lo = {f_5,f_4,f_3,f_2,f_1,1'h0}; // @[Cat.scala 31:58]
  wire [11:0] io_f_lo_lo = {f_11,f_10,f_9,f_8,f_7,f_6,io_f_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] io_f_lo_hi_lo = {f_17,f_16,f_15,f_14,f_13,f_12}; // @[Cat.scala 31:58]
  wire [23:0] io_f_lo = {f_23,f_22,f_21,f_20,f_19,f_18,io_f_lo_hi_lo,io_f_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] io_f_hi_lo_lo = {f_29,f_28,f_27,f_26,f_25,f_24}; // @[Cat.scala 31:58]
  wire [11:0] io_f_hi_lo = {f_35,f_34,f_33,f_32,f_31,f_30,io_f_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] io_f_hi_hi_lo = {f_41,f_40,f_39,f_38,f_37,f_36}; // @[Cat.scala 31:58]
  wire [24:0] io_f_hi = {f_48,f_47,f_46,f_45,f_44,f_43,f_42,io_f_hi_hi_lo,io_f_hi_lo}; // @[Cat.scala 31:58]
  assign io_f = {io_f_hi,io_f_lo}; // @[Cat.scala 31:58]
endmodule

